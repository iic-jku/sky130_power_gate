magic
tech sky130A
magscale 1 2
timestamp 1697797845
<< locali >>
rect 36 22768 1802 22958
rect 36 21986 340 22768
rect 870 21986 1802 22768
rect 36 21800 1802 21986
<< viali >>
rect 340 21986 870 22768
<< metal1 >>
rect 122 45072 132 45126
rect 1706 45072 1716 45126
rect 132 682 178 45072
rect 1660 23168 1706 45072
rect 334 22768 876 22780
rect 330 21986 340 22768
rect 870 21986 880 22768
rect 334 21974 876 21986
rect 1660 632 1708 23168
rect 1660 584 1706 632
<< via1 >>
rect 132 45072 1706 45126
rect 340 21986 870 22768
<< metal2 >>
rect 132 45136 1706 45146
rect 132 45052 1706 45062
rect 340 22768 870 22778
rect 340 21976 870 21986
<< via2 >>
rect 132 45126 1706 45136
rect 132 45072 1706 45126
rect 132 45062 1706 45072
rect 340 21986 870 22768
<< metal3 >>
rect 122 45136 1716 45141
rect 122 45062 132 45136
rect 1706 45062 1716 45136
rect 122 45057 1716 45062
rect 330 22768 880 22773
rect 330 21986 340 22768
rect 870 21986 880 22768
rect 330 21981 880 21986
<< via3 >>
rect 132 45062 1706 45136
rect 340 21986 870 22768
<< metal4 >>
rect 0 45136 1840 45152
rect 0 45062 132 45136
rect 1706 45062 1840 45136
rect 0 45052 1840 45062
rect 0 0 240 44848
rect 340 22769 870 44848
rect 339 22768 871 22769
rect 339 21986 340 22768
rect 870 21986 871 22768
rect 339 21985 871 21986
rect 340 0 870 21985
rect 970 0 1500 44848
rect 1600 0 1840 44848
use pmos  pmos_0
timestamp 1697796922
transform 1 0 0 0 1 22408
box 0 490 1838 21944
use pmos  pmos_1
timestamp 1697796922
transform 1 0 0 0 1 -90
box 0 490 1838 21944
<< labels >>
rlabel metal4 0 0 240 44848 1 VGND
port 1 n ground input
rlabel metal4 1600 0 1840 44848 1 VGND
port 1 n ground input
rlabel metal4 340 0 870 44848 1 VPWR
port 2 n power input
rlabel metal4 970 0 1500 44848 1 GPWR
port 3 n power output
rlabel metal4 0 45052 1840 45152 1 ctrl
port 4 n signal input
<< end >>
