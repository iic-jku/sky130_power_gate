magic
tech sky130A
magscale 1 2
timestamp 1685958313
<< locali >>
rect -1370 692 -1356 696
rect -1370 -292 -1252 692
rect -1326 -720 -1252 -292
rect -1370 -914 -1252 -720
rect -756 -916 -638 694
<< viali >>
rect -934 836 11098 872
rect -1390 -720 -1326 -292
<< metal1 >>
rect -946 872 11110 878
rect -946 830 -934 872
rect -944 814 -934 830
rect 11098 830 11110 872
rect -708 810 -702 814
rect 11098 810 11108 830
rect -1244 752 -762 776
rect -1244 722 -744 752
rect -650 730 10980 778
rect -1178 238 -836 690
rect -1178 220 -834 238
rect -1168 20 -834 220
rect -780 78 -770 690
rect -708 78 -698 690
rect -650 20 -602 730
rect -464 90 -454 690
rect -396 90 -386 690
rect -272 90 -262 690
rect -204 90 -194 690
rect -80 90 -70 690
rect -12 90 -2 690
rect 112 90 122 690
rect 180 90 190 690
rect 304 90 314 690
rect 372 90 382 690
rect 496 90 506 690
rect 564 90 574 690
rect 688 90 698 690
rect 756 90 766 690
rect 880 90 890 690
rect 948 90 958 690
rect 1072 90 1082 690
rect 1140 90 1150 690
rect 1264 88 1274 688
rect 1332 88 1342 688
rect 1456 88 1466 688
rect 1524 88 1534 688
rect 1648 88 1658 688
rect 1716 88 1726 688
rect 1840 88 1850 688
rect 1908 88 1918 688
rect 2032 88 2042 688
rect 2100 88 2110 688
rect 2224 88 2234 688
rect 2292 88 2302 688
rect 2416 88 2426 688
rect 2484 88 2494 688
rect 2608 88 2618 688
rect 2676 88 2686 688
rect 2800 88 2810 688
rect 2868 88 2878 688
rect 2992 88 3002 688
rect 3060 88 3070 688
rect 3184 88 3194 688
rect 3252 88 3262 688
rect 3376 88 3386 688
rect 3444 88 3454 688
rect 3568 88 3578 688
rect 3636 88 3646 688
rect 3760 88 3770 688
rect 3828 88 3838 688
rect 3952 88 3962 688
rect 4020 88 4030 688
rect 4144 88 4154 688
rect 4212 88 4222 688
rect 4336 88 4346 688
rect 4404 88 4414 688
rect 4528 88 4538 688
rect 4596 88 4606 688
rect 4720 88 4730 688
rect 4788 88 4798 688
rect 4912 88 4922 688
rect 4980 88 4990 688
rect 5104 88 5114 688
rect 5172 88 5182 688
rect 5296 88 5306 688
rect 5364 88 5374 688
rect 5488 88 5498 688
rect 5556 88 5566 688
rect 5680 88 5690 688
rect 5748 88 5758 688
rect 5872 88 5882 688
rect 5940 88 5950 688
rect 6064 88 6074 688
rect 6132 88 6142 688
rect 6256 88 6266 688
rect 6324 88 6334 688
rect 6448 88 6458 688
rect 6516 88 6526 688
rect 6640 88 6650 688
rect 6708 88 6718 688
rect 6832 88 6842 688
rect 6900 88 6910 688
rect 7024 88 7034 688
rect 7092 88 7102 688
rect 7216 88 7226 688
rect 7284 88 7294 688
rect 7408 88 7418 688
rect 7476 88 7486 688
rect 7600 88 7610 688
rect 7668 88 7678 688
rect 7792 88 7802 688
rect 7860 88 7870 688
rect 7984 88 7994 688
rect 8052 88 8062 688
rect 8176 88 8186 688
rect 8244 88 8254 688
rect 8368 88 8378 688
rect 8436 88 8446 688
rect 8560 88 8570 688
rect 8628 88 8638 688
rect 8752 88 8762 688
rect 8820 88 8830 688
rect 8944 88 8954 688
rect 9012 88 9022 688
rect 9136 88 9146 688
rect 9204 88 9214 688
rect 9328 88 9338 688
rect 9396 88 9406 688
rect 9520 88 9530 688
rect 9588 88 9598 688
rect 9712 88 9722 688
rect 9780 88 9790 688
rect 9904 88 9914 688
rect 9972 88 9982 688
rect 10096 88 10106 688
rect 10164 88 10174 688
rect 10288 88 10298 688
rect 10356 88 10366 688
rect 10480 88 10490 688
rect 10548 88 10558 688
rect 10672 88 10682 688
rect 10740 88 10750 688
rect 10864 88 10874 688
rect 10932 88 10942 688
rect -1168 -52 -978 20
rect -1172 -80 -978 -52
rect -1178 -228 -978 -80
rect -896 -94 -834 20
rect -896 -228 -836 -94
rect -694 -228 -684 20
rect -602 -228 -592 20
rect -1400 -292 -1272 -280
rect -1400 -720 -1390 -292
rect -1326 -668 -1272 -292
rect -1326 -720 -1258 -668
rect -1400 -732 -1258 -720
rect -1178 -910 -836 -228
rect -1256 -1000 -1246 -942
rect -1094 -1000 -764 -942
rect -650 -952 -602 -228
rect -560 -912 -550 -312
rect -492 -912 -482 -312
rect -368 -912 -358 -312
rect -300 -912 -290 -312
rect -176 -912 -166 -312
rect -108 -912 -98 -312
rect 16 -912 26 -312
rect 84 -912 94 -312
rect 208 -912 218 -312
rect 276 -912 286 -312
rect 400 -912 410 -312
rect 468 -912 478 -312
rect 592 -912 602 -312
rect 660 -912 670 -312
rect 784 -912 794 -312
rect 852 -912 862 -312
rect 976 -912 986 -312
rect 1044 -912 1054 -312
rect 1168 -912 1178 -312
rect 1236 -912 1246 -312
rect 1360 -912 1370 -312
rect 1428 -912 1438 -312
rect 1552 -912 1562 -312
rect 1620 -912 1630 -312
rect 1744 -912 1754 -312
rect 1812 -912 1822 -312
rect 1936 -912 1946 -312
rect 2004 -912 2014 -312
rect 2128 -912 2138 -312
rect 2196 -912 2206 -312
rect 2320 -912 2330 -312
rect 2388 -912 2398 -312
rect 2512 -912 2522 -312
rect 2580 -912 2590 -312
rect 2704 -912 2714 -312
rect 2772 -912 2782 -312
rect 2896 -912 2906 -312
rect 2964 -912 2974 -312
rect 3088 -912 3098 -312
rect 3156 -912 3166 -312
rect 3280 -912 3290 -312
rect 3348 -912 3358 -312
rect 3472 -912 3482 -312
rect 3540 -912 3550 -312
rect 3664 -912 3674 -312
rect 3732 -912 3742 -312
rect 3856 -912 3866 -312
rect 3924 -912 3934 -312
rect 4048 -912 4058 -312
rect 4116 -912 4126 -312
rect 4240 -912 4250 -312
rect 4308 -912 4318 -312
rect 4432 -912 4442 -312
rect 4500 -912 4510 -312
rect 4624 -912 4634 -312
rect 4692 -912 4702 -312
rect 4816 -912 4826 -312
rect 4884 -912 4894 -312
rect 5008 -912 5018 -312
rect 5076 -912 5086 -312
rect 5200 -912 5210 -312
rect 5268 -912 5278 -312
rect 5392 -912 5402 -312
rect 5460 -912 5470 -312
rect 5584 -912 5594 -312
rect 5652 -912 5662 -312
rect 5776 -912 5786 -312
rect 5844 -912 5854 -312
rect 5968 -912 5978 -312
rect 6036 -912 6046 -312
rect 6160 -912 6170 -312
rect 6228 -912 6238 -312
rect 6352 -912 6362 -312
rect 6420 -912 6430 -312
rect 6544 -912 6554 -312
rect 6612 -912 6622 -312
rect 6736 -912 6746 -312
rect 6804 -912 6814 -312
rect 6928 -912 6938 -312
rect 6996 -912 7006 -312
rect 7120 -912 7130 -312
rect 7188 -912 7198 -312
rect 7312 -912 7322 -312
rect 7380 -912 7390 -312
rect 7504 -912 7514 -312
rect 7572 -912 7582 -312
rect 7696 -912 7706 -312
rect 7764 -912 7774 -312
rect 7888 -912 7898 -312
rect 7956 -912 7966 -312
rect 8080 -912 8090 -312
rect 8148 -912 8158 -312
rect 8272 -912 8282 -312
rect 8340 -912 8350 -312
rect 8464 -912 8474 -312
rect 8532 -912 8542 -312
rect 8656 -912 8666 -312
rect 8724 -912 8734 -312
rect 8848 -912 8858 -312
rect 8916 -912 8926 -312
rect 9040 -912 9050 -312
rect 9108 -912 9118 -312
rect 9232 -912 9242 -312
rect 9300 -912 9310 -312
rect 9424 -912 9434 -312
rect 9492 -912 9502 -312
rect 9616 -912 9626 -312
rect 9684 -912 9694 -312
rect 9808 -912 9818 -312
rect 9876 -912 9886 -312
rect 10000 -912 10010 -312
rect 10068 -912 10078 -312
rect 10192 -912 10202 -312
rect 10260 -912 10270 -312
rect 10384 -912 10394 -312
rect 10452 -912 10462 -312
rect 10576 -912 10586 -312
rect 10644 -912 10654 -312
rect 10768 -912 10778 -312
rect 10836 -912 10846 -312
rect 10960 -912 10970 -312
rect 11028 -912 11038 -312
rect -650 -1000 10884 -952
<< via1 >>
rect -934 836 11098 872
rect -934 814 11098 836
rect -702 810 11098 814
rect -770 78 -708 690
rect -454 90 -396 690
rect -262 90 -204 690
rect -70 90 -12 690
rect 122 90 180 690
rect 314 90 372 690
rect 506 90 564 690
rect 698 90 756 690
rect 890 90 948 690
rect 1082 90 1140 690
rect 1274 88 1332 688
rect 1466 88 1524 688
rect 1658 88 1716 688
rect 1850 88 1908 688
rect 2042 88 2100 688
rect 2234 88 2292 688
rect 2426 88 2484 688
rect 2618 88 2676 688
rect 2810 88 2868 688
rect 3002 88 3060 688
rect 3194 88 3252 688
rect 3386 88 3444 688
rect 3578 88 3636 688
rect 3770 88 3828 688
rect 3962 88 4020 688
rect 4154 88 4212 688
rect 4346 88 4404 688
rect 4538 88 4596 688
rect 4730 88 4788 688
rect 4922 88 4980 688
rect 5114 88 5172 688
rect 5306 88 5364 688
rect 5498 88 5556 688
rect 5690 88 5748 688
rect 5882 88 5940 688
rect 6074 88 6132 688
rect 6266 88 6324 688
rect 6458 88 6516 688
rect 6650 88 6708 688
rect 6842 88 6900 688
rect 7034 88 7092 688
rect 7226 88 7284 688
rect 7418 88 7476 688
rect 7610 88 7668 688
rect 7802 88 7860 688
rect 7994 88 8052 688
rect 8186 88 8244 688
rect 8378 88 8436 688
rect 8570 88 8628 688
rect 8762 88 8820 688
rect 8954 88 9012 688
rect 9146 88 9204 688
rect 9338 88 9396 688
rect 9530 88 9588 688
rect 9722 88 9780 688
rect 9914 88 9972 688
rect 10106 88 10164 688
rect 10298 88 10356 688
rect 10490 88 10548 688
rect 10682 88 10740 688
rect 10874 88 10932 688
rect -978 -228 -896 20
rect -684 -228 -602 20
rect -1390 -720 -1326 -292
rect -1246 -1000 -1094 -942
rect -550 -912 -492 -312
rect -358 -912 -300 -312
rect -166 -912 -108 -312
rect 26 -912 84 -312
rect 218 -912 276 -312
rect 410 -912 468 -312
rect 602 -912 660 -312
rect 794 -912 852 -312
rect 986 -912 1044 -312
rect 1178 -912 1236 -312
rect 1370 -912 1428 -312
rect 1562 -912 1620 -312
rect 1754 -912 1812 -312
rect 1946 -912 2004 -312
rect 2138 -912 2196 -312
rect 2330 -912 2388 -312
rect 2522 -912 2580 -312
rect 2714 -912 2772 -312
rect 2906 -912 2964 -312
rect 3098 -912 3156 -312
rect 3290 -912 3348 -312
rect 3482 -912 3540 -312
rect 3674 -912 3732 -312
rect 3866 -912 3924 -312
rect 4058 -912 4116 -312
rect 4250 -912 4308 -312
rect 4442 -912 4500 -312
rect 4634 -912 4692 -312
rect 4826 -912 4884 -312
rect 5018 -912 5076 -312
rect 5210 -912 5268 -312
rect 5402 -912 5460 -312
rect 5594 -912 5652 -312
rect 5786 -912 5844 -312
rect 5978 -912 6036 -312
rect 6170 -912 6228 -312
rect 6362 -912 6420 -312
rect 6554 -912 6612 -312
rect 6746 -912 6804 -312
rect 6938 -912 6996 -312
rect 7130 -912 7188 -312
rect 7322 -912 7380 -312
rect 7514 -912 7572 -312
rect 7706 -912 7764 -312
rect 7898 -912 7956 -312
rect 8090 -912 8148 -312
rect 8282 -912 8340 -312
rect 8474 -912 8532 -312
rect 8666 -912 8724 -312
rect 8858 -912 8916 -312
rect 9050 -912 9108 -312
rect 9242 -912 9300 -312
rect 9434 -912 9492 -312
rect 9626 -912 9684 -312
rect 9818 -912 9876 -312
rect 10010 -912 10068 -312
rect 10202 -912 10260 -312
rect 10394 -912 10452 -312
rect 10586 -912 10644 -312
rect 10778 -912 10836 -312
rect 10970 -912 11028 -312
<< metal2 >>
rect -934 872 11098 882
rect -934 800 11098 810
rect -770 690 -708 800
rect -770 68 -708 78
rect -454 698 10934 708
rect -454 70 10934 80
rect -978 20 -602 32
rect -896 -228 -684 20
rect -978 -238 -602 -228
rect -1390 -292 -1326 -282
rect -1390 -730 -1326 -720
rect -550 -302 11028 -292
rect -1416 -922 -1094 -912
rect -550 -932 11028 -922
rect -1416 -1030 -1094 -1020
<< via2 >>
rect -934 814 11098 872
rect -934 810 -702 814
rect -702 810 11098 814
rect -454 690 10934 698
rect -454 90 -396 690
rect -396 90 -262 690
rect -262 90 -204 690
rect -204 90 -70 690
rect -70 90 -12 690
rect -12 90 122 690
rect 122 90 180 690
rect 180 90 314 690
rect 314 90 372 690
rect 372 90 506 690
rect 506 90 564 690
rect 564 90 698 690
rect 698 90 756 690
rect 756 90 890 690
rect 890 90 948 690
rect 948 90 1082 690
rect 1082 90 1140 690
rect 1140 688 10934 690
rect 1140 90 1274 688
rect -454 88 1274 90
rect 1274 88 1332 688
rect 1332 88 1466 688
rect 1466 88 1524 688
rect 1524 88 1658 688
rect 1658 88 1716 688
rect 1716 88 1850 688
rect 1850 88 1908 688
rect 1908 88 2042 688
rect 2042 88 2100 688
rect 2100 88 2234 688
rect 2234 88 2292 688
rect 2292 88 2426 688
rect 2426 88 2484 688
rect 2484 88 2618 688
rect 2618 88 2676 688
rect 2676 88 2810 688
rect 2810 88 2868 688
rect 2868 88 3002 688
rect 3002 88 3060 688
rect 3060 88 3194 688
rect 3194 88 3252 688
rect 3252 88 3386 688
rect 3386 88 3444 688
rect 3444 88 3578 688
rect 3578 88 3636 688
rect 3636 88 3770 688
rect 3770 88 3828 688
rect 3828 88 3962 688
rect 3962 88 4020 688
rect 4020 88 4154 688
rect 4154 88 4212 688
rect 4212 88 4346 688
rect 4346 88 4404 688
rect 4404 88 4538 688
rect 4538 88 4596 688
rect 4596 88 4730 688
rect 4730 88 4788 688
rect 4788 88 4922 688
rect 4922 88 4980 688
rect 4980 88 5114 688
rect 5114 88 5172 688
rect 5172 88 5306 688
rect 5306 88 5364 688
rect 5364 88 5498 688
rect 5498 88 5556 688
rect 5556 88 5690 688
rect 5690 88 5748 688
rect 5748 88 5882 688
rect 5882 88 5940 688
rect 5940 88 6074 688
rect 6074 88 6132 688
rect 6132 88 6266 688
rect 6266 88 6324 688
rect 6324 88 6458 688
rect 6458 88 6516 688
rect 6516 88 6650 688
rect 6650 88 6708 688
rect 6708 88 6842 688
rect 6842 88 6900 688
rect 6900 88 7034 688
rect 7034 88 7092 688
rect 7092 88 7226 688
rect 7226 88 7284 688
rect 7284 88 7418 688
rect 7418 88 7476 688
rect 7476 88 7610 688
rect 7610 88 7668 688
rect 7668 88 7802 688
rect 7802 88 7860 688
rect 7860 88 7994 688
rect 7994 88 8052 688
rect 8052 88 8186 688
rect 8186 88 8244 688
rect 8244 88 8378 688
rect 8378 88 8436 688
rect 8436 88 8570 688
rect 8570 88 8628 688
rect 8628 88 8762 688
rect 8762 88 8820 688
rect 8820 88 8954 688
rect 8954 88 9012 688
rect 9012 88 9146 688
rect 9146 88 9204 688
rect 9204 88 9338 688
rect 9338 88 9396 688
rect 9396 88 9530 688
rect 9530 88 9588 688
rect 9588 88 9722 688
rect 9722 88 9780 688
rect 9780 88 9914 688
rect 9914 88 9972 688
rect 9972 88 10106 688
rect 10106 88 10164 688
rect 10164 88 10298 688
rect 10298 88 10356 688
rect 10356 88 10490 688
rect 10490 88 10548 688
rect 10548 88 10682 688
rect 10682 88 10740 688
rect 10740 88 10874 688
rect 10874 88 10932 688
rect 10932 88 10934 688
rect -454 80 10934 88
rect -1390 -720 -1326 -292
rect -550 -312 11028 -302
rect -550 -912 -492 -312
rect -492 -912 -358 -312
rect -358 -912 -300 -312
rect -300 -912 -166 -312
rect -166 -912 -108 -312
rect -108 -912 26 -312
rect 26 -912 84 -312
rect 84 -912 218 -312
rect 218 -912 276 -312
rect 276 -912 410 -312
rect 410 -912 468 -312
rect 468 -912 602 -312
rect 602 -912 660 -312
rect 660 -912 794 -312
rect 794 -912 852 -312
rect 852 -912 986 -312
rect 986 -912 1044 -312
rect 1044 -912 1178 -312
rect 1178 -912 1236 -312
rect 1236 -912 1370 -312
rect 1370 -912 1428 -312
rect 1428 -912 1562 -312
rect 1562 -912 1620 -312
rect 1620 -912 1754 -312
rect 1754 -912 1812 -312
rect 1812 -912 1946 -312
rect 1946 -912 2004 -312
rect 2004 -912 2138 -312
rect 2138 -912 2196 -312
rect 2196 -912 2330 -312
rect 2330 -912 2388 -312
rect 2388 -912 2522 -312
rect 2522 -912 2580 -312
rect 2580 -912 2714 -312
rect 2714 -912 2772 -312
rect 2772 -912 2906 -312
rect 2906 -912 2964 -312
rect 2964 -912 3098 -312
rect 3098 -912 3156 -312
rect 3156 -912 3290 -312
rect 3290 -912 3348 -312
rect 3348 -912 3482 -312
rect 3482 -912 3540 -312
rect 3540 -912 3674 -312
rect 3674 -912 3732 -312
rect 3732 -912 3866 -312
rect 3866 -912 3924 -312
rect 3924 -912 4058 -312
rect 4058 -912 4116 -312
rect 4116 -912 4250 -312
rect 4250 -912 4308 -312
rect 4308 -912 4442 -312
rect 4442 -912 4500 -312
rect 4500 -912 4634 -312
rect 4634 -912 4692 -312
rect 4692 -912 4826 -312
rect 4826 -912 4884 -312
rect 4884 -912 5018 -312
rect 5018 -912 5076 -312
rect 5076 -912 5210 -312
rect 5210 -912 5268 -312
rect 5268 -912 5402 -312
rect 5402 -912 5460 -312
rect 5460 -912 5594 -312
rect 5594 -912 5652 -312
rect 5652 -912 5786 -312
rect 5786 -912 5844 -312
rect 5844 -912 5978 -312
rect 5978 -912 6036 -312
rect 6036 -912 6170 -312
rect 6170 -912 6228 -312
rect 6228 -912 6362 -312
rect 6362 -912 6420 -312
rect 6420 -912 6554 -312
rect 6554 -912 6612 -312
rect 6612 -912 6746 -312
rect 6746 -912 6804 -312
rect 6804 -912 6938 -312
rect 6938 -912 6996 -312
rect 6996 -912 7130 -312
rect 7130 -912 7188 -312
rect 7188 -912 7322 -312
rect 7322 -912 7380 -312
rect 7380 -912 7514 -312
rect 7514 -912 7572 -312
rect 7572 -912 7706 -312
rect 7706 -912 7764 -312
rect 7764 -912 7898 -312
rect 7898 -912 7956 -312
rect 7956 -912 8090 -312
rect 8090 -912 8148 -312
rect 8148 -912 8282 -312
rect 8282 -912 8340 -312
rect 8340 -912 8474 -312
rect 8474 -912 8532 -312
rect 8532 -912 8666 -312
rect 8666 -912 8724 -312
rect 8724 -912 8858 -312
rect 8858 -912 8916 -312
rect 8916 -912 9050 -312
rect 9050 -912 9108 -312
rect 9108 -912 9242 -312
rect 9242 -912 9300 -312
rect 9300 -912 9434 -312
rect 9434 -912 9492 -312
rect 9492 -912 9626 -312
rect 9626 -912 9684 -312
rect 9684 -912 9818 -312
rect 9818 -912 9876 -312
rect 9876 -912 10010 -312
rect 10010 -912 10068 -312
rect 10068 -912 10202 -312
rect 10202 -912 10260 -312
rect 10260 -912 10394 -312
rect 10394 -912 10452 -312
rect 10452 -912 10586 -312
rect 10586 -912 10644 -312
rect 10644 -912 10778 -312
rect 10778 -912 10836 -312
rect 10836 -912 10970 -312
rect 10970 -912 11028 -312
rect -1416 -942 -1094 -922
rect -550 -922 11028 -912
rect -1416 -1000 -1246 -942
rect -1246 -1000 -1094 -942
rect -1416 -1020 -1094 -1000
<< metal3 >>
rect -1428 872 11166 908
rect -1428 810 -934 872
rect 11098 810 11166 872
rect -1428 698 11166 810
rect -1428 80 -454 698
rect 10934 80 11166 698
rect -464 75 11166 80
rect 10934 74 11166 75
rect -1400 -292 -1316 -287
rect -1426 -720 -1390 -292
rect -1326 -720 -1088 -292
rect -1426 -722 -1088 -720
rect -1006 -302 11168 -292
rect -1400 -725 -1316 -722
rect -1426 -922 -1088 -916
rect -1426 -1020 -1416 -922
rect -1094 -1020 -1088 -922
rect -1426 -1134 -1088 -1020
rect -1006 -922 -550 -302
rect 11028 -922 11168 -302
rect -1006 -1134 11168 -922
use sky130_fd_pr__nfet_01v8_H2P3K4  sky130_fd_pr__nfet_01v8_H2P3K4_0
timestamp 1685732482
transform 1 0 -1215 0 1 -110
box -210 -1010 210 1010
use sky130_fd_pr__pfet_01v8_3QZTZS  sky130_fd_pr__pfet_01v8_3QZTZS_0
timestamp 1685741491
transform 1 0 5239 0 1 -111
box -5926 -1018 5926 1018
use sky130_fd_pr__pfet_01v8_XYJ9AL  sky130_fd_pr__pfet_01v8_XYJ9AL_0
timestamp 1685740367
transform 1 0 -791 0 1 -111
box -210 -1018 210 1018
<< labels >>
rlabel metal3 -1428 698 11166 908 1 vdd
port 1 n default bidirectional
rlabel metal3 -1006 -1134 11168 -922 1 vdd_switch
port 4 n default bidirectional
rlabel metal3 -1426 -722 -1088 -292 1 vss
port 3 n default bidirectional
rlabel metal3 -1426 -1134 -1088 -916 1 en
port 2 n default input
<< end >>
