magic
tech sky130A
magscale 1 2
timestamp 1697193306
<< nwell >>
rect 0 546 1838 22000
<< pmos >>
rect 219 21770 1619 21800
rect 219 21674 1619 21704
rect 219 21578 1619 21608
rect 219 21482 1619 21512
rect 219 21386 1619 21416
rect 219 21290 1619 21320
rect 219 21194 1619 21224
rect 219 21098 1619 21128
rect 219 21002 1619 21032
rect 219 20906 1619 20936
rect 219 20810 1619 20840
rect 219 20714 1619 20744
rect 219 20618 1619 20648
rect 219 20522 1619 20552
rect 219 20426 1619 20456
rect 219 20330 1619 20360
rect 219 20234 1619 20264
rect 219 20138 1619 20168
rect 219 20042 1619 20072
rect 219 19946 1619 19976
rect 219 19850 1619 19880
rect 219 19754 1619 19784
rect 219 19658 1619 19688
rect 219 19562 1619 19592
rect 219 19466 1619 19496
rect 219 19370 1619 19400
rect 219 19274 1619 19304
rect 219 19178 1619 19208
rect 219 19082 1619 19112
rect 219 18986 1619 19016
rect 219 18890 1619 18920
rect 219 18794 1619 18824
rect 219 18698 1619 18728
rect 219 18602 1619 18632
rect 219 18506 1619 18536
rect 219 18410 1619 18440
rect 219 18314 1619 18344
rect 219 18218 1619 18248
rect 219 18122 1619 18152
rect 219 18026 1619 18056
rect 219 17930 1619 17960
rect 219 17834 1619 17864
rect 219 17738 1619 17768
rect 219 17642 1619 17672
rect 219 17546 1619 17576
rect 219 17450 1619 17480
rect 219 17354 1619 17384
rect 219 17258 1619 17288
rect 219 17162 1619 17192
rect 219 17066 1619 17096
rect 219 16970 1619 17000
rect 219 16874 1619 16904
rect 219 16778 1619 16808
rect 219 16682 1619 16712
rect 219 16586 1619 16616
rect 219 16490 1619 16520
rect 219 16394 1619 16424
rect 219 16298 1619 16328
rect 219 16202 1619 16232
rect 219 16106 1619 16136
rect 219 16010 1619 16040
rect 219 15914 1619 15944
rect 219 15818 1619 15848
rect 219 15722 1619 15752
rect 219 15626 1619 15656
rect 219 15530 1619 15560
rect 219 15434 1619 15464
rect 219 15338 1619 15368
rect 219 15242 1619 15272
rect 219 15146 1619 15176
rect 219 15050 1619 15080
rect 219 14954 1619 14984
rect 219 14858 1619 14888
rect 219 14762 1619 14792
rect 219 14666 1619 14696
rect 219 14570 1619 14600
rect 219 14474 1619 14504
rect 219 14378 1619 14408
rect 219 14282 1619 14312
rect 219 14186 1619 14216
rect 219 14090 1619 14120
rect 219 13994 1619 14024
rect 219 13898 1619 13928
rect 219 13802 1619 13832
rect 219 13706 1619 13736
rect 219 13610 1619 13640
rect 219 13514 1619 13544
rect 219 13418 1619 13448
rect 219 13322 1619 13352
rect 219 13226 1619 13256
rect 219 13130 1619 13160
rect 219 13034 1619 13064
rect 219 12938 1619 12968
rect 219 12842 1619 12872
rect 219 12746 1619 12776
rect 219 12650 1619 12680
rect 219 12554 1619 12584
rect 219 12458 1619 12488
rect 219 12362 1619 12392
rect 219 12266 1619 12296
rect 219 12170 1619 12200
rect 219 12074 1619 12104
rect 219 11978 1619 12008
rect 219 11882 1619 11912
rect 219 11786 1619 11816
rect 219 11690 1619 11720
rect 219 11594 1619 11624
rect 219 11498 1619 11528
rect 219 11402 1619 11432
rect 219 11306 1619 11336
rect 219 11210 1619 11240
rect 219 11114 1619 11144
rect 219 11018 1619 11048
rect 219 10922 1619 10952
rect 219 10826 1619 10856
rect 219 10730 1619 10760
rect 219 10634 1619 10664
rect 219 10538 1619 10568
rect 219 10442 1619 10472
rect 219 10346 1619 10376
rect 219 10250 1619 10280
rect 219 10154 1619 10184
rect 219 10058 1619 10088
rect 219 9962 1619 9992
rect 219 9866 1619 9896
rect 219 9770 1619 9800
rect 219 9674 1619 9704
rect 219 9578 1619 9608
rect 219 9482 1619 9512
rect 219 9386 1619 9416
rect 219 9290 1619 9320
rect 219 9194 1619 9224
rect 219 9098 1619 9128
rect 219 9002 1619 9032
rect 219 8906 1619 8936
rect 219 8810 1619 8840
rect 219 8714 1619 8744
rect 219 8618 1619 8648
rect 219 8522 1619 8552
rect 219 8426 1619 8456
rect 219 8330 1619 8360
rect 219 8234 1619 8264
rect 219 8138 1619 8168
rect 219 8042 1619 8072
rect 219 7946 1619 7976
rect 219 7850 1619 7880
rect 219 7754 1619 7784
rect 219 7658 1619 7688
rect 219 7562 1619 7592
rect 219 7466 1619 7496
rect 219 7370 1619 7400
rect 219 7274 1619 7304
rect 219 7178 1619 7208
rect 219 7082 1619 7112
rect 219 6986 1619 7016
rect 219 6890 1619 6920
rect 219 6794 1619 6824
rect 219 6698 1619 6728
rect 219 6602 1619 6632
rect 219 6506 1619 6536
rect 219 6410 1619 6440
rect 219 6314 1619 6344
rect 219 6218 1619 6248
rect 219 6122 1619 6152
rect 219 6026 1619 6056
rect 219 5930 1619 5960
rect 219 5834 1619 5864
rect 219 5738 1619 5768
rect 219 5642 1619 5672
rect 219 5546 1619 5576
rect 219 5450 1619 5480
rect 219 5354 1619 5384
rect 219 5258 1619 5288
rect 219 5162 1619 5192
rect 219 5066 1619 5096
rect 219 4970 1619 5000
rect 219 4874 1619 4904
rect 219 4778 1619 4808
rect 219 4682 1619 4712
rect 219 4586 1619 4616
rect 219 4490 1619 4520
rect 219 4394 1619 4424
rect 219 4298 1619 4328
rect 219 4202 1619 4232
rect 219 4106 1619 4136
rect 219 4010 1619 4040
rect 219 3914 1619 3944
rect 219 3818 1619 3848
rect 219 3722 1619 3752
rect 219 3626 1619 3656
rect 219 3530 1619 3560
rect 219 3434 1619 3464
rect 219 3338 1619 3368
rect 219 3242 1619 3272
rect 219 3146 1619 3176
rect 219 3050 1619 3080
rect 219 2954 1619 2984
rect 219 2858 1619 2888
rect 219 2762 1619 2792
rect 219 2666 1619 2696
rect 219 2570 1619 2600
rect 219 2474 1619 2504
rect 219 2378 1619 2408
rect 219 2282 1619 2312
rect 219 2186 1619 2216
rect 219 2090 1619 2120
rect 219 1994 1619 2024
rect 219 1898 1619 1928
rect 219 1802 1619 1832
rect 219 1706 1619 1736
rect 219 1610 1619 1640
rect 219 1514 1619 1544
rect 219 1418 1619 1448
rect 219 1322 1619 1352
rect 219 1226 1619 1256
rect 219 1130 1619 1160
rect 219 1034 1619 1064
rect 219 938 1619 968
rect 219 842 1619 872
rect 219 746 1619 776
<< pdiff >>
rect 219 21850 1619 21862
rect 219 21816 231 21850
rect 1607 21816 1619 21850
rect 219 21800 1619 21816
rect 219 21754 1619 21770
rect 219 21720 231 21754
rect 1607 21720 1619 21754
rect 219 21704 1619 21720
rect 219 21658 1619 21674
rect 219 21624 231 21658
rect 1607 21624 1619 21658
rect 219 21608 1619 21624
rect 219 21562 1619 21578
rect 219 21528 231 21562
rect 1607 21528 1619 21562
rect 219 21512 1619 21528
rect 219 21466 1619 21482
rect 219 21432 231 21466
rect 1607 21432 1619 21466
rect 219 21416 1619 21432
rect 219 21370 1619 21386
rect 219 21336 231 21370
rect 1607 21336 1619 21370
rect 219 21320 1619 21336
rect 219 21274 1619 21290
rect 219 21240 231 21274
rect 1607 21240 1619 21274
rect 219 21224 1619 21240
rect 219 21178 1619 21194
rect 219 21144 231 21178
rect 1607 21144 1619 21178
rect 219 21128 1619 21144
rect 219 21082 1619 21098
rect 219 21048 231 21082
rect 1607 21048 1619 21082
rect 219 21032 1619 21048
rect 219 20986 1619 21002
rect 219 20952 231 20986
rect 1607 20952 1619 20986
rect 219 20936 1619 20952
rect 219 20890 1619 20906
rect 219 20856 231 20890
rect 1607 20856 1619 20890
rect 219 20840 1619 20856
rect 219 20794 1619 20810
rect 219 20760 231 20794
rect 1607 20760 1619 20794
rect 219 20744 1619 20760
rect 219 20698 1619 20714
rect 219 20664 231 20698
rect 1607 20664 1619 20698
rect 219 20648 1619 20664
rect 219 20602 1619 20618
rect 219 20568 231 20602
rect 1607 20568 1619 20602
rect 219 20552 1619 20568
rect 219 20506 1619 20522
rect 219 20472 231 20506
rect 1607 20472 1619 20506
rect 219 20456 1619 20472
rect 219 20410 1619 20426
rect 219 20376 231 20410
rect 1607 20376 1619 20410
rect 219 20360 1619 20376
rect 219 20314 1619 20330
rect 219 20280 231 20314
rect 1607 20280 1619 20314
rect 219 20264 1619 20280
rect 219 20218 1619 20234
rect 219 20184 231 20218
rect 1607 20184 1619 20218
rect 219 20168 1619 20184
rect 219 20122 1619 20138
rect 219 20088 231 20122
rect 1607 20088 1619 20122
rect 219 20072 1619 20088
rect 219 20026 1619 20042
rect 219 19992 231 20026
rect 1607 19992 1619 20026
rect 219 19976 1619 19992
rect 219 19930 1619 19946
rect 219 19896 231 19930
rect 1607 19896 1619 19930
rect 219 19880 1619 19896
rect 219 19834 1619 19850
rect 219 19800 231 19834
rect 1607 19800 1619 19834
rect 219 19784 1619 19800
rect 219 19738 1619 19754
rect 219 19704 231 19738
rect 1607 19704 1619 19738
rect 219 19688 1619 19704
rect 219 19642 1619 19658
rect 219 19608 231 19642
rect 1607 19608 1619 19642
rect 219 19592 1619 19608
rect 219 19546 1619 19562
rect 219 19512 231 19546
rect 1607 19512 1619 19546
rect 219 19496 1619 19512
rect 219 19450 1619 19466
rect 219 19416 231 19450
rect 1607 19416 1619 19450
rect 219 19400 1619 19416
rect 219 19354 1619 19370
rect 219 19320 231 19354
rect 1607 19320 1619 19354
rect 219 19304 1619 19320
rect 219 19258 1619 19274
rect 219 19224 231 19258
rect 1607 19224 1619 19258
rect 219 19208 1619 19224
rect 219 19162 1619 19178
rect 219 19128 231 19162
rect 1607 19128 1619 19162
rect 219 19112 1619 19128
rect 219 19066 1619 19082
rect 219 19032 231 19066
rect 1607 19032 1619 19066
rect 219 19016 1619 19032
rect 219 18970 1619 18986
rect 219 18936 231 18970
rect 1607 18936 1619 18970
rect 219 18920 1619 18936
rect 219 18874 1619 18890
rect 219 18840 231 18874
rect 1607 18840 1619 18874
rect 219 18824 1619 18840
rect 219 18778 1619 18794
rect 219 18744 231 18778
rect 1607 18744 1619 18778
rect 219 18728 1619 18744
rect 219 18682 1619 18698
rect 219 18648 231 18682
rect 1607 18648 1619 18682
rect 219 18632 1619 18648
rect 219 18586 1619 18602
rect 219 18552 231 18586
rect 1607 18552 1619 18586
rect 219 18536 1619 18552
rect 219 18490 1619 18506
rect 219 18456 231 18490
rect 1607 18456 1619 18490
rect 219 18440 1619 18456
rect 219 18394 1619 18410
rect 219 18360 231 18394
rect 1607 18360 1619 18394
rect 219 18344 1619 18360
rect 219 18298 1619 18314
rect 219 18264 231 18298
rect 1607 18264 1619 18298
rect 219 18248 1619 18264
rect 219 18202 1619 18218
rect 219 18168 231 18202
rect 1607 18168 1619 18202
rect 219 18152 1619 18168
rect 219 18106 1619 18122
rect 219 18072 231 18106
rect 1607 18072 1619 18106
rect 219 18056 1619 18072
rect 219 18010 1619 18026
rect 219 17976 231 18010
rect 1607 17976 1619 18010
rect 219 17960 1619 17976
rect 219 17914 1619 17930
rect 219 17880 231 17914
rect 1607 17880 1619 17914
rect 219 17864 1619 17880
rect 219 17818 1619 17834
rect 219 17784 231 17818
rect 1607 17784 1619 17818
rect 219 17768 1619 17784
rect 219 17722 1619 17738
rect 219 17688 231 17722
rect 1607 17688 1619 17722
rect 219 17672 1619 17688
rect 219 17626 1619 17642
rect 219 17592 231 17626
rect 1607 17592 1619 17626
rect 219 17576 1619 17592
rect 219 17530 1619 17546
rect 219 17496 231 17530
rect 1607 17496 1619 17530
rect 219 17480 1619 17496
rect 219 17434 1619 17450
rect 219 17400 231 17434
rect 1607 17400 1619 17434
rect 219 17384 1619 17400
rect 219 17338 1619 17354
rect 219 17304 231 17338
rect 1607 17304 1619 17338
rect 219 17288 1619 17304
rect 219 17242 1619 17258
rect 219 17208 231 17242
rect 1607 17208 1619 17242
rect 219 17192 1619 17208
rect 219 17146 1619 17162
rect 219 17112 231 17146
rect 1607 17112 1619 17146
rect 219 17096 1619 17112
rect 219 17050 1619 17066
rect 219 17016 231 17050
rect 1607 17016 1619 17050
rect 219 17000 1619 17016
rect 219 16954 1619 16970
rect 219 16920 231 16954
rect 1607 16920 1619 16954
rect 219 16904 1619 16920
rect 219 16858 1619 16874
rect 219 16824 231 16858
rect 1607 16824 1619 16858
rect 219 16808 1619 16824
rect 219 16762 1619 16778
rect 219 16728 231 16762
rect 1607 16728 1619 16762
rect 219 16712 1619 16728
rect 219 16666 1619 16682
rect 219 16632 231 16666
rect 1607 16632 1619 16666
rect 219 16616 1619 16632
rect 219 16570 1619 16586
rect 219 16536 231 16570
rect 1607 16536 1619 16570
rect 219 16520 1619 16536
rect 219 16474 1619 16490
rect 219 16440 231 16474
rect 1607 16440 1619 16474
rect 219 16424 1619 16440
rect 219 16378 1619 16394
rect 219 16344 231 16378
rect 1607 16344 1619 16378
rect 219 16328 1619 16344
rect 219 16282 1619 16298
rect 219 16248 231 16282
rect 1607 16248 1619 16282
rect 219 16232 1619 16248
rect 219 16186 1619 16202
rect 219 16152 231 16186
rect 1607 16152 1619 16186
rect 219 16136 1619 16152
rect 219 16090 1619 16106
rect 219 16056 231 16090
rect 1607 16056 1619 16090
rect 219 16040 1619 16056
rect 219 15994 1619 16010
rect 219 15960 231 15994
rect 1607 15960 1619 15994
rect 219 15944 1619 15960
rect 219 15898 1619 15914
rect 219 15864 231 15898
rect 1607 15864 1619 15898
rect 219 15848 1619 15864
rect 219 15802 1619 15818
rect 219 15768 231 15802
rect 1607 15768 1619 15802
rect 219 15752 1619 15768
rect 219 15706 1619 15722
rect 219 15672 231 15706
rect 1607 15672 1619 15706
rect 219 15656 1619 15672
rect 219 15610 1619 15626
rect 219 15576 231 15610
rect 1607 15576 1619 15610
rect 219 15560 1619 15576
rect 219 15514 1619 15530
rect 219 15480 231 15514
rect 1607 15480 1619 15514
rect 219 15464 1619 15480
rect 219 15418 1619 15434
rect 219 15384 231 15418
rect 1607 15384 1619 15418
rect 219 15368 1619 15384
rect 219 15322 1619 15338
rect 219 15288 231 15322
rect 1607 15288 1619 15322
rect 219 15272 1619 15288
rect 219 15226 1619 15242
rect 219 15192 231 15226
rect 1607 15192 1619 15226
rect 219 15176 1619 15192
rect 219 15130 1619 15146
rect 219 15096 231 15130
rect 1607 15096 1619 15130
rect 219 15080 1619 15096
rect 219 15034 1619 15050
rect 219 15000 231 15034
rect 1607 15000 1619 15034
rect 219 14984 1619 15000
rect 219 14938 1619 14954
rect 219 14904 231 14938
rect 1607 14904 1619 14938
rect 219 14888 1619 14904
rect 219 14842 1619 14858
rect 219 14808 231 14842
rect 1607 14808 1619 14842
rect 219 14792 1619 14808
rect 219 14746 1619 14762
rect 219 14712 231 14746
rect 1607 14712 1619 14746
rect 219 14696 1619 14712
rect 219 14650 1619 14666
rect 219 14616 231 14650
rect 1607 14616 1619 14650
rect 219 14600 1619 14616
rect 219 14554 1619 14570
rect 219 14520 231 14554
rect 1607 14520 1619 14554
rect 219 14504 1619 14520
rect 219 14458 1619 14474
rect 219 14424 231 14458
rect 1607 14424 1619 14458
rect 219 14408 1619 14424
rect 219 14362 1619 14378
rect 219 14328 231 14362
rect 1607 14328 1619 14362
rect 219 14312 1619 14328
rect 219 14266 1619 14282
rect 219 14232 231 14266
rect 1607 14232 1619 14266
rect 219 14216 1619 14232
rect 219 14170 1619 14186
rect 219 14136 231 14170
rect 1607 14136 1619 14170
rect 219 14120 1619 14136
rect 219 14074 1619 14090
rect 219 14040 231 14074
rect 1607 14040 1619 14074
rect 219 14024 1619 14040
rect 219 13978 1619 13994
rect 219 13944 231 13978
rect 1607 13944 1619 13978
rect 219 13928 1619 13944
rect 219 13882 1619 13898
rect 219 13848 231 13882
rect 1607 13848 1619 13882
rect 219 13832 1619 13848
rect 219 13786 1619 13802
rect 219 13752 231 13786
rect 1607 13752 1619 13786
rect 219 13736 1619 13752
rect 219 13690 1619 13706
rect 219 13656 231 13690
rect 1607 13656 1619 13690
rect 219 13640 1619 13656
rect 219 13594 1619 13610
rect 219 13560 231 13594
rect 1607 13560 1619 13594
rect 219 13544 1619 13560
rect 219 13498 1619 13514
rect 219 13464 231 13498
rect 1607 13464 1619 13498
rect 219 13448 1619 13464
rect 219 13402 1619 13418
rect 219 13368 231 13402
rect 1607 13368 1619 13402
rect 219 13352 1619 13368
rect 219 13306 1619 13322
rect 219 13272 231 13306
rect 1607 13272 1619 13306
rect 219 13256 1619 13272
rect 219 13210 1619 13226
rect 219 13176 231 13210
rect 1607 13176 1619 13210
rect 219 13160 1619 13176
rect 219 13114 1619 13130
rect 219 13080 231 13114
rect 1607 13080 1619 13114
rect 219 13064 1619 13080
rect 219 13018 1619 13034
rect 219 12984 231 13018
rect 1607 12984 1619 13018
rect 219 12968 1619 12984
rect 219 12922 1619 12938
rect 219 12888 231 12922
rect 1607 12888 1619 12922
rect 219 12872 1619 12888
rect 219 12826 1619 12842
rect 219 12792 231 12826
rect 1607 12792 1619 12826
rect 219 12776 1619 12792
rect 219 12730 1619 12746
rect 219 12696 231 12730
rect 1607 12696 1619 12730
rect 219 12680 1619 12696
rect 219 12634 1619 12650
rect 219 12600 231 12634
rect 1607 12600 1619 12634
rect 219 12584 1619 12600
rect 219 12538 1619 12554
rect 219 12504 231 12538
rect 1607 12504 1619 12538
rect 219 12488 1619 12504
rect 219 12442 1619 12458
rect 219 12408 231 12442
rect 1607 12408 1619 12442
rect 219 12392 1619 12408
rect 219 12346 1619 12362
rect 219 12312 231 12346
rect 1607 12312 1619 12346
rect 219 12296 1619 12312
rect 219 12250 1619 12266
rect 219 12216 231 12250
rect 1607 12216 1619 12250
rect 219 12200 1619 12216
rect 219 12154 1619 12170
rect 219 12120 231 12154
rect 1607 12120 1619 12154
rect 219 12104 1619 12120
rect 219 12058 1619 12074
rect 219 12024 231 12058
rect 1607 12024 1619 12058
rect 219 12008 1619 12024
rect 219 11962 1619 11978
rect 219 11928 231 11962
rect 1607 11928 1619 11962
rect 219 11912 1619 11928
rect 219 11866 1619 11882
rect 219 11832 231 11866
rect 1607 11832 1619 11866
rect 219 11816 1619 11832
rect 219 11770 1619 11786
rect 219 11736 231 11770
rect 1607 11736 1619 11770
rect 219 11720 1619 11736
rect 219 11674 1619 11690
rect 219 11640 231 11674
rect 1607 11640 1619 11674
rect 219 11624 1619 11640
rect 219 11578 1619 11594
rect 219 11544 231 11578
rect 1607 11544 1619 11578
rect 219 11528 1619 11544
rect 219 11482 1619 11498
rect 219 11448 231 11482
rect 1607 11448 1619 11482
rect 219 11432 1619 11448
rect 219 11386 1619 11402
rect 219 11352 231 11386
rect 1607 11352 1619 11386
rect 219 11336 1619 11352
rect 219 11290 1619 11306
rect 219 11256 231 11290
rect 1607 11256 1619 11290
rect 219 11240 1619 11256
rect 219 11194 1619 11210
rect 219 11160 231 11194
rect 1607 11160 1619 11194
rect 219 11144 1619 11160
rect 219 11098 1619 11114
rect 219 11064 231 11098
rect 1607 11064 1619 11098
rect 219 11048 1619 11064
rect 219 11002 1619 11018
rect 219 10968 231 11002
rect 1607 10968 1619 11002
rect 219 10952 1619 10968
rect 219 10906 1619 10922
rect 219 10872 231 10906
rect 1607 10872 1619 10906
rect 219 10856 1619 10872
rect 219 10810 1619 10826
rect 219 10776 231 10810
rect 1607 10776 1619 10810
rect 219 10760 1619 10776
rect 219 10714 1619 10730
rect 219 10680 231 10714
rect 1607 10680 1619 10714
rect 219 10664 1619 10680
rect 219 10618 1619 10634
rect 219 10584 231 10618
rect 1607 10584 1619 10618
rect 219 10568 1619 10584
rect 219 10522 1619 10538
rect 219 10488 231 10522
rect 1607 10488 1619 10522
rect 219 10472 1619 10488
rect 219 10426 1619 10442
rect 219 10392 231 10426
rect 1607 10392 1619 10426
rect 219 10376 1619 10392
rect 219 10330 1619 10346
rect 219 10296 231 10330
rect 1607 10296 1619 10330
rect 219 10280 1619 10296
rect 219 10234 1619 10250
rect 219 10200 231 10234
rect 1607 10200 1619 10234
rect 219 10184 1619 10200
rect 219 10138 1619 10154
rect 219 10104 231 10138
rect 1607 10104 1619 10138
rect 219 10088 1619 10104
rect 219 10042 1619 10058
rect 219 10008 231 10042
rect 1607 10008 1619 10042
rect 219 9992 1619 10008
rect 219 9946 1619 9962
rect 219 9912 231 9946
rect 1607 9912 1619 9946
rect 219 9896 1619 9912
rect 219 9850 1619 9866
rect 219 9816 231 9850
rect 1607 9816 1619 9850
rect 219 9800 1619 9816
rect 219 9754 1619 9770
rect 219 9720 231 9754
rect 1607 9720 1619 9754
rect 219 9704 1619 9720
rect 219 9658 1619 9674
rect 219 9624 231 9658
rect 1607 9624 1619 9658
rect 219 9608 1619 9624
rect 219 9562 1619 9578
rect 219 9528 231 9562
rect 1607 9528 1619 9562
rect 219 9512 1619 9528
rect 219 9466 1619 9482
rect 219 9432 231 9466
rect 1607 9432 1619 9466
rect 219 9416 1619 9432
rect 219 9370 1619 9386
rect 219 9336 231 9370
rect 1607 9336 1619 9370
rect 219 9320 1619 9336
rect 219 9274 1619 9290
rect 219 9240 231 9274
rect 1607 9240 1619 9274
rect 219 9224 1619 9240
rect 219 9178 1619 9194
rect 219 9144 231 9178
rect 1607 9144 1619 9178
rect 219 9128 1619 9144
rect 219 9082 1619 9098
rect 219 9048 231 9082
rect 1607 9048 1619 9082
rect 219 9032 1619 9048
rect 219 8986 1619 9002
rect 219 8952 231 8986
rect 1607 8952 1619 8986
rect 219 8936 1619 8952
rect 219 8890 1619 8906
rect 219 8856 231 8890
rect 1607 8856 1619 8890
rect 219 8840 1619 8856
rect 219 8794 1619 8810
rect 219 8760 231 8794
rect 1607 8760 1619 8794
rect 219 8744 1619 8760
rect 219 8698 1619 8714
rect 219 8664 231 8698
rect 1607 8664 1619 8698
rect 219 8648 1619 8664
rect 219 8602 1619 8618
rect 219 8568 231 8602
rect 1607 8568 1619 8602
rect 219 8552 1619 8568
rect 219 8506 1619 8522
rect 219 8472 231 8506
rect 1607 8472 1619 8506
rect 219 8456 1619 8472
rect 219 8410 1619 8426
rect 219 8376 231 8410
rect 1607 8376 1619 8410
rect 219 8360 1619 8376
rect 219 8314 1619 8330
rect 219 8280 231 8314
rect 1607 8280 1619 8314
rect 219 8264 1619 8280
rect 219 8218 1619 8234
rect 219 8184 231 8218
rect 1607 8184 1619 8218
rect 219 8168 1619 8184
rect 219 8122 1619 8138
rect 219 8088 231 8122
rect 1607 8088 1619 8122
rect 219 8072 1619 8088
rect 219 8026 1619 8042
rect 219 7992 231 8026
rect 1607 7992 1619 8026
rect 219 7976 1619 7992
rect 219 7930 1619 7946
rect 219 7896 231 7930
rect 1607 7896 1619 7930
rect 219 7880 1619 7896
rect 219 7834 1619 7850
rect 219 7800 231 7834
rect 1607 7800 1619 7834
rect 219 7784 1619 7800
rect 219 7738 1619 7754
rect 219 7704 231 7738
rect 1607 7704 1619 7738
rect 219 7688 1619 7704
rect 219 7642 1619 7658
rect 219 7608 231 7642
rect 1607 7608 1619 7642
rect 219 7592 1619 7608
rect 219 7546 1619 7562
rect 219 7512 231 7546
rect 1607 7512 1619 7546
rect 219 7496 1619 7512
rect 219 7450 1619 7466
rect 219 7416 231 7450
rect 1607 7416 1619 7450
rect 219 7400 1619 7416
rect 219 7354 1619 7370
rect 219 7320 231 7354
rect 1607 7320 1619 7354
rect 219 7304 1619 7320
rect 219 7258 1619 7274
rect 219 7224 231 7258
rect 1607 7224 1619 7258
rect 219 7208 1619 7224
rect 219 7162 1619 7178
rect 219 7128 231 7162
rect 1607 7128 1619 7162
rect 219 7112 1619 7128
rect 219 7066 1619 7082
rect 219 7032 231 7066
rect 1607 7032 1619 7066
rect 219 7016 1619 7032
rect 219 6970 1619 6986
rect 219 6936 231 6970
rect 1607 6936 1619 6970
rect 219 6920 1619 6936
rect 219 6874 1619 6890
rect 219 6840 231 6874
rect 1607 6840 1619 6874
rect 219 6824 1619 6840
rect 219 6778 1619 6794
rect 219 6744 231 6778
rect 1607 6744 1619 6778
rect 219 6728 1619 6744
rect 219 6682 1619 6698
rect 219 6648 231 6682
rect 1607 6648 1619 6682
rect 219 6632 1619 6648
rect 219 6586 1619 6602
rect 219 6552 231 6586
rect 1607 6552 1619 6586
rect 219 6536 1619 6552
rect 219 6490 1619 6506
rect 219 6456 231 6490
rect 1607 6456 1619 6490
rect 219 6440 1619 6456
rect 219 6394 1619 6410
rect 219 6360 231 6394
rect 1607 6360 1619 6394
rect 219 6344 1619 6360
rect 219 6298 1619 6314
rect 219 6264 231 6298
rect 1607 6264 1619 6298
rect 219 6248 1619 6264
rect 219 6202 1619 6218
rect 219 6168 231 6202
rect 1607 6168 1619 6202
rect 219 6152 1619 6168
rect 219 6106 1619 6122
rect 219 6072 231 6106
rect 1607 6072 1619 6106
rect 219 6056 1619 6072
rect 219 6010 1619 6026
rect 219 5976 231 6010
rect 1607 5976 1619 6010
rect 219 5960 1619 5976
rect 219 5914 1619 5930
rect 219 5880 231 5914
rect 1607 5880 1619 5914
rect 219 5864 1619 5880
rect 219 5818 1619 5834
rect 219 5784 231 5818
rect 1607 5784 1619 5818
rect 219 5768 1619 5784
rect 219 5722 1619 5738
rect 219 5688 231 5722
rect 1607 5688 1619 5722
rect 219 5672 1619 5688
rect 219 5626 1619 5642
rect 219 5592 231 5626
rect 1607 5592 1619 5626
rect 219 5576 1619 5592
rect 219 5530 1619 5546
rect 219 5496 231 5530
rect 1607 5496 1619 5530
rect 219 5480 1619 5496
rect 219 5434 1619 5450
rect 219 5400 231 5434
rect 1607 5400 1619 5434
rect 219 5384 1619 5400
rect 219 5338 1619 5354
rect 219 5304 231 5338
rect 1607 5304 1619 5338
rect 219 5288 1619 5304
rect 219 5242 1619 5258
rect 219 5208 231 5242
rect 1607 5208 1619 5242
rect 219 5192 1619 5208
rect 219 5146 1619 5162
rect 219 5112 231 5146
rect 1607 5112 1619 5146
rect 219 5096 1619 5112
rect 219 5050 1619 5066
rect 219 5016 231 5050
rect 1607 5016 1619 5050
rect 219 5000 1619 5016
rect 219 4954 1619 4970
rect 219 4920 231 4954
rect 1607 4920 1619 4954
rect 219 4904 1619 4920
rect 219 4858 1619 4874
rect 219 4824 231 4858
rect 1607 4824 1619 4858
rect 219 4808 1619 4824
rect 219 4762 1619 4778
rect 219 4728 231 4762
rect 1607 4728 1619 4762
rect 219 4712 1619 4728
rect 219 4666 1619 4682
rect 219 4632 231 4666
rect 1607 4632 1619 4666
rect 219 4616 1619 4632
rect 219 4570 1619 4586
rect 219 4536 231 4570
rect 1607 4536 1619 4570
rect 219 4520 1619 4536
rect 219 4474 1619 4490
rect 219 4440 231 4474
rect 1607 4440 1619 4474
rect 219 4424 1619 4440
rect 219 4378 1619 4394
rect 219 4344 231 4378
rect 1607 4344 1619 4378
rect 219 4328 1619 4344
rect 219 4282 1619 4298
rect 219 4248 231 4282
rect 1607 4248 1619 4282
rect 219 4232 1619 4248
rect 219 4186 1619 4202
rect 219 4152 231 4186
rect 1607 4152 1619 4186
rect 219 4136 1619 4152
rect 219 4090 1619 4106
rect 219 4056 231 4090
rect 1607 4056 1619 4090
rect 219 4040 1619 4056
rect 219 3994 1619 4010
rect 219 3960 231 3994
rect 1607 3960 1619 3994
rect 219 3944 1619 3960
rect 219 3898 1619 3914
rect 219 3864 231 3898
rect 1607 3864 1619 3898
rect 219 3848 1619 3864
rect 219 3802 1619 3818
rect 219 3768 231 3802
rect 1607 3768 1619 3802
rect 219 3752 1619 3768
rect 219 3706 1619 3722
rect 219 3672 231 3706
rect 1607 3672 1619 3706
rect 219 3656 1619 3672
rect 219 3610 1619 3626
rect 219 3576 231 3610
rect 1607 3576 1619 3610
rect 219 3560 1619 3576
rect 219 3514 1619 3530
rect 219 3480 231 3514
rect 1607 3480 1619 3514
rect 219 3464 1619 3480
rect 219 3418 1619 3434
rect 219 3384 231 3418
rect 1607 3384 1619 3418
rect 219 3368 1619 3384
rect 219 3322 1619 3338
rect 219 3288 231 3322
rect 1607 3288 1619 3322
rect 219 3272 1619 3288
rect 219 3226 1619 3242
rect 219 3192 231 3226
rect 1607 3192 1619 3226
rect 219 3176 1619 3192
rect 219 3130 1619 3146
rect 219 3096 231 3130
rect 1607 3096 1619 3130
rect 219 3080 1619 3096
rect 219 3034 1619 3050
rect 219 3000 231 3034
rect 1607 3000 1619 3034
rect 219 2984 1619 3000
rect 219 2938 1619 2954
rect 219 2904 231 2938
rect 1607 2904 1619 2938
rect 219 2888 1619 2904
rect 219 2842 1619 2858
rect 219 2808 231 2842
rect 1607 2808 1619 2842
rect 219 2792 1619 2808
rect 219 2746 1619 2762
rect 219 2712 231 2746
rect 1607 2712 1619 2746
rect 219 2696 1619 2712
rect 219 2650 1619 2666
rect 219 2616 231 2650
rect 1607 2616 1619 2650
rect 219 2600 1619 2616
rect 219 2554 1619 2570
rect 219 2520 231 2554
rect 1607 2520 1619 2554
rect 219 2504 1619 2520
rect 219 2458 1619 2474
rect 219 2424 231 2458
rect 1607 2424 1619 2458
rect 219 2408 1619 2424
rect 219 2362 1619 2378
rect 219 2328 231 2362
rect 1607 2328 1619 2362
rect 219 2312 1619 2328
rect 219 2266 1619 2282
rect 219 2232 231 2266
rect 1607 2232 1619 2266
rect 219 2216 1619 2232
rect 219 2170 1619 2186
rect 219 2136 231 2170
rect 1607 2136 1619 2170
rect 219 2120 1619 2136
rect 219 2074 1619 2090
rect 219 2040 231 2074
rect 1607 2040 1619 2074
rect 219 2024 1619 2040
rect 219 1978 1619 1994
rect 219 1944 231 1978
rect 1607 1944 1619 1978
rect 219 1928 1619 1944
rect 219 1882 1619 1898
rect 219 1848 231 1882
rect 1607 1848 1619 1882
rect 219 1832 1619 1848
rect 219 1786 1619 1802
rect 219 1752 231 1786
rect 1607 1752 1619 1786
rect 219 1736 1619 1752
rect 219 1690 1619 1706
rect 219 1656 231 1690
rect 1607 1656 1619 1690
rect 219 1640 1619 1656
rect 219 1594 1619 1610
rect 219 1560 231 1594
rect 1607 1560 1619 1594
rect 219 1544 1619 1560
rect 219 1498 1619 1514
rect 219 1464 231 1498
rect 1607 1464 1619 1498
rect 219 1448 1619 1464
rect 219 1402 1619 1418
rect 219 1368 231 1402
rect 1607 1368 1619 1402
rect 219 1352 1619 1368
rect 219 1306 1619 1322
rect 219 1272 231 1306
rect 1607 1272 1619 1306
rect 219 1256 1619 1272
rect 219 1210 1619 1226
rect 219 1176 231 1210
rect 1607 1176 1619 1210
rect 219 1160 1619 1176
rect 219 1114 1619 1130
rect 219 1080 231 1114
rect 1607 1080 1619 1114
rect 219 1064 1619 1080
rect 219 1018 1619 1034
rect 219 984 231 1018
rect 1607 984 1619 1018
rect 219 968 1619 984
rect 219 922 1619 938
rect 219 888 231 922
rect 1607 888 1619 922
rect 219 872 1619 888
rect 219 826 1619 842
rect 219 792 231 826
rect 1607 792 1619 826
rect 219 776 1619 792
rect 219 730 1619 746
rect 219 696 231 730
rect 1607 696 1619 730
rect 219 684 1619 696
<< pdiffc >>
rect 231 21816 1607 21850
rect 231 21720 1607 21754
rect 231 21624 1607 21658
rect 231 21528 1607 21562
rect 231 21432 1607 21466
rect 231 21336 1607 21370
rect 231 21240 1607 21274
rect 231 21144 1607 21178
rect 231 21048 1607 21082
rect 231 20952 1607 20986
rect 231 20856 1607 20890
rect 231 20760 1607 20794
rect 231 20664 1607 20698
rect 231 20568 1607 20602
rect 231 20472 1607 20506
rect 231 20376 1607 20410
rect 231 20280 1607 20314
rect 231 20184 1607 20218
rect 231 20088 1607 20122
rect 231 19992 1607 20026
rect 231 19896 1607 19930
rect 231 19800 1607 19834
rect 231 19704 1607 19738
rect 231 19608 1607 19642
rect 231 19512 1607 19546
rect 231 19416 1607 19450
rect 231 19320 1607 19354
rect 231 19224 1607 19258
rect 231 19128 1607 19162
rect 231 19032 1607 19066
rect 231 18936 1607 18970
rect 231 18840 1607 18874
rect 231 18744 1607 18778
rect 231 18648 1607 18682
rect 231 18552 1607 18586
rect 231 18456 1607 18490
rect 231 18360 1607 18394
rect 231 18264 1607 18298
rect 231 18168 1607 18202
rect 231 18072 1607 18106
rect 231 17976 1607 18010
rect 231 17880 1607 17914
rect 231 17784 1607 17818
rect 231 17688 1607 17722
rect 231 17592 1607 17626
rect 231 17496 1607 17530
rect 231 17400 1607 17434
rect 231 17304 1607 17338
rect 231 17208 1607 17242
rect 231 17112 1607 17146
rect 231 17016 1607 17050
rect 231 16920 1607 16954
rect 231 16824 1607 16858
rect 231 16728 1607 16762
rect 231 16632 1607 16666
rect 231 16536 1607 16570
rect 231 16440 1607 16474
rect 231 16344 1607 16378
rect 231 16248 1607 16282
rect 231 16152 1607 16186
rect 231 16056 1607 16090
rect 231 15960 1607 15994
rect 231 15864 1607 15898
rect 231 15768 1607 15802
rect 231 15672 1607 15706
rect 231 15576 1607 15610
rect 231 15480 1607 15514
rect 231 15384 1607 15418
rect 231 15288 1607 15322
rect 231 15192 1607 15226
rect 231 15096 1607 15130
rect 231 15000 1607 15034
rect 231 14904 1607 14938
rect 231 14808 1607 14842
rect 231 14712 1607 14746
rect 231 14616 1607 14650
rect 231 14520 1607 14554
rect 231 14424 1607 14458
rect 231 14328 1607 14362
rect 231 14232 1607 14266
rect 231 14136 1607 14170
rect 231 14040 1607 14074
rect 231 13944 1607 13978
rect 231 13848 1607 13882
rect 231 13752 1607 13786
rect 231 13656 1607 13690
rect 231 13560 1607 13594
rect 231 13464 1607 13498
rect 231 13368 1607 13402
rect 231 13272 1607 13306
rect 231 13176 1607 13210
rect 231 13080 1607 13114
rect 231 12984 1607 13018
rect 231 12888 1607 12922
rect 231 12792 1607 12826
rect 231 12696 1607 12730
rect 231 12600 1607 12634
rect 231 12504 1607 12538
rect 231 12408 1607 12442
rect 231 12312 1607 12346
rect 231 12216 1607 12250
rect 231 12120 1607 12154
rect 231 12024 1607 12058
rect 231 11928 1607 11962
rect 231 11832 1607 11866
rect 231 11736 1607 11770
rect 231 11640 1607 11674
rect 231 11544 1607 11578
rect 231 11448 1607 11482
rect 231 11352 1607 11386
rect 231 11256 1607 11290
rect 231 11160 1607 11194
rect 231 11064 1607 11098
rect 231 10968 1607 11002
rect 231 10872 1607 10906
rect 231 10776 1607 10810
rect 231 10680 1607 10714
rect 231 10584 1607 10618
rect 231 10488 1607 10522
rect 231 10392 1607 10426
rect 231 10296 1607 10330
rect 231 10200 1607 10234
rect 231 10104 1607 10138
rect 231 10008 1607 10042
rect 231 9912 1607 9946
rect 231 9816 1607 9850
rect 231 9720 1607 9754
rect 231 9624 1607 9658
rect 231 9528 1607 9562
rect 231 9432 1607 9466
rect 231 9336 1607 9370
rect 231 9240 1607 9274
rect 231 9144 1607 9178
rect 231 9048 1607 9082
rect 231 8952 1607 8986
rect 231 8856 1607 8890
rect 231 8760 1607 8794
rect 231 8664 1607 8698
rect 231 8568 1607 8602
rect 231 8472 1607 8506
rect 231 8376 1607 8410
rect 231 8280 1607 8314
rect 231 8184 1607 8218
rect 231 8088 1607 8122
rect 231 7992 1607 8026
rect 231 7896 1607 7930
rect 231 7800 1607 7834
rect 231 7704 1607 7738
rect 231 7608 1607 7642
rect 231 7512 1607 7546
rect 231 7416 1607 7450
rect 231 7320 1607 7354
rect 231 7224 1607 7258
rect 231 7128 1607 7162
rect 231 7032 1607 7066
rect 231 6936 1607 6970
rect 231 6840 1607 6874
rect 231 6744 1607 6778
rect 231 6648 1607 6682
rect 231 6552 1607 6586
rect 231 6456 1607 6490
rect 231 6360 1607 6394
rect 231 6264 1607 6298
rect 231 6168 1607 6202
rect 231 6072 1607 6106
rect 231 5976 1607 6010
rect 231 5880 1607 5914
rect 231 5784 1607 5818
rect 231 5688 1607 5722
rect 231 5592 1607 5626
rect 231 5496 1607 5530
rect 231 5400 1607 5434
rect 231 5304 1607 5338
rect 231 5208 1607 5242
rect 231 5112 1607 5146
rect 231 5016 1607 5050
rect 231 4920 1607 4954
rect 231 4824 1607 4858
rect 231 4728 1607 4762
rect 231 4632 1607 4666
rect 231 4536 1607 4570
rect 231 4440 1607 4474
rect 231 4344 1607 4378
rect 231 4248 1607 4282
rect 231 4152 1607 4186
rect 231 4056 1607 4090
rect 231 3960 1607 3994
rect 231 3864 1607 3898
rect 231 3768 1607 3802
rect 231 3672 1607 3706
rect 231 3576 1607 3610
rect 231 3480 1607 3514
rect 231 3384 1607 3418
rect 231 3288 1607 3322
rect 231 3192 1607 3226
rect 231 3096 1607 3130
rect 231 3000 1607 3034
rect 231 2904 1607 2938
rect 231 2808 1607 2842
rect 231 2712 1607 2746
rect 231 2616 1607 2650
rect 231 2520 1607 2554
rect 231 2424 1607 2458
rect 231 2328 1607 2362
rect 231 2232 1607 2266
rect 231 2136 1607 2170
rect 231 2040 1607 2074
rect 231 1944 1607 1978
rect 231 1848 1607 1882
rect 231 1752 1607 1786
rect 231 1656 1607 1690
rect 231 1560 1607 1594
rect 231 1464 1607 1498
rect 231 1368 1607 1402
rect 231 1272 1607 1306
rect 231 1176 1607 1210
rect 231 1080 1607 1114
rect 231 984 1607 1018
rect 231 888 1607 922
rect 231 792 1607 826
rect 231 696 1607 730
<< nsubdiff >>
rect 36 21930 132 21964
rect 1706 21930 1802 21964
rect 36 21868 70 21930
rect 1768 21868 1802 21930
rect 36 616 70 678
rect 1768 616 1802 678
rect 36 582 132 616
rect 1706 582 1802 616
<< nsubdiffcont >>
rect 132 21930 1706 21964
rect 36 678 70 21868
rect 1768 678 1802 21868
rect 132 582 1706 616
<< poly >>
rect 122 21802 188 21818
rect 122 21768 138 21802
rect 172 21800 188 21802
rect 172 21770 219 21800
rect 1619 21770 1645 21800
rect 172 21768 188 21770
rect 122 21752 188 21768
rect 1650 21706 1716 21722
rect 1650 21704 1666 21706
rect 193 21674 219 21704
rect 1619 21674 1666 21704
rect 122 21610 188 21626
rect 122 21576 138 21610
rect 172 21608 188 21610
rect 1650 21672 1666 21674
rect 1700 21672 1716 21706
rect 1650 21656 1716 21672
rect 172 21578 219 21608
rect 1619 21578 1645 21608
rect 172 21576 188 21578
rect 122 21560 188 21576
rect 1650 21514 1716 21530
rect 1650 21512 1666 21514
rect 193 21482 219 21512
rect 1619 21482 1666 21512
rect 122 21418 188 21434
rect 122 21384 138 21418
rect 172 21416 188 21418
rect 1650 21480 1666 21482
rect 1700 21480 1716 21514
rect 1650 21464 1716 21480
rect 172 21386 219 21416
rect 1619 21386 1645 21416
rect 172 21384 188 21386
rect 122 21368 188 21384
rect 1650 21322 1716 21338
rect 1650 21320 1666 21322
rect 193 21290 219 21320
rect 1619 21290 1666 21320
rect 122 21226 188 21242
rect 122 21192 138 21226
rect 172 21224 188 21226
rect 1650 21288 1666 21290
rect 1700 21288 1716 21322
rect 1650 21272 1716 21288
rect 172 21194 219 21224
rect 1619 21194 1645 21224
rect 172 21192 188 21194
rect 122 21176 188 21192
rect 1650 21130 1716 21146
rect 1650 21128 1666 21130
rect 193 21098 219 21128
rect 1619 21098 1666 21128
rect 122 21034 188 21050
rect 122 21000 138 21034
rect 172 21032 188 21034
rect 1650 21096 1666 21098
rect 1700 21096 1716 21130
rect 1650 21080 1716 21096
rect 172 21002 219 21032
rect 1619 21002 1645 21032
rect 172 21000 188 21002
rect 122 20984 188 21000
rect 1650 20938 1716 20954
rect 1650 20936 1666 20938
rect 193 20906 219 20936
rect 1619 20906 1666 20936
rect 122 20842 188 20858
rect 122 20808 138 20842
rect 172 20840 188 20842
rect 1650 20904 1666 20906
rect 1700 20904 1716 20938
rect 1650 20888 1716 20904
rect 172 20810 219 20840
rect 1619 20810 1645 20840
rect 172 20808 188 20810
rect 122 20792 188 20808
rect 1650 20746 1716 20762
rect 1650 20744 1666 20746
rect 193 20714 219 20744
rect 1619 20714 1666 20744
rect 122 20650 188 20666
rect 122 20616 138 20650
rect 172 20648 188 20650
rect 1650 20712 1666 20714
rect 1700 20712 1716 20746
rect 1650 20696 1716 20712
rect 172 20618 219 20648
rect 1619 20618 1645 20648
rect 172 20616 188 20618
rect 122 20600 188 20616
rect 1650 20554 1716 20570
rect 1650 20552 1666 20554
rect 193 20522 219 20552
rect 1619 20522 1666 20552
rect 122 20458 188 20474
rect 122 20424 138 20458
rect 172 20456 188 20458
rect 1650 20520 1666 20522
rect 1700 20520 1716 20554
rect 1650 20504 1716 20520
rect 172 20426 219 20456
rect 1619 20426 1645 20456
rect 172 20424 188 20426
rect 122 20408 188 20424
rect 1650 20362 1716 20378
rect 1650 20360 1666 20362
rect 193 20330 219 20360
rect 1619 20330 1666 20360
rect 122 20266 188 20282
rect 122 20232 138 20266
rect 172 20264 188 20266
rect 1650 20328 1666 20330
rect 1700 20328 1716 20362
rect 1650 20312 1716 20328
rect 172 20234 219 20264
rect 1619 20234 1645 20264
rect 172 20232 188 20234
rect 122 20216 188 20232
rect 1650 20170 1716 20186
rect 1650 20168 1666 20170
rect 193 20138 219 20168
rect 1619 20138 1666 20168
rect 122 20074 188 20090
rect 122 20040 138 20074
rect 172 20072 188 20074
rect 1650 20136 1666 20138
rect 1700 20136 1716 20170
rect 1650 20120 1716 20136
rect 172 20042 219 20072
rect 1619 20042 1645 20072
rect 172 20040 188 20042
rect 122 20024 188 20040
rect 1650 19978 1716 19994
rect 1650 19976 1666 19978
rect 193 19946 219 19976
rect 1619 19946 1666 19976
rect 122 19882 188 19898
rect 122 19848 138 19882
rect 172 19880 188 19882
rect 1650 19944 1666 19946
rect 1700 19944 1716 19978
rect 1650 19928 1716 19944
rect 172 19850 219 19880
rect 1619 19850 1645 19880
rect 172 19848 188 19850
rect 122 19832 188 19848
rect 1650 19786 1716 19802
rect 1650 19784 1666 19786
rect 193 19754 219 19784
rect 1619 19754 1666 19784
rect 122 19690 188 19706
rect 122 19656 138 19690
rect 172 19688 188 19690
rect 1650 19752 1666 19754
rect 1700 19752 1716 19786
rect 1650 19736 1716 19752
rect 172 19658 219 19688
rect 1619 19658 1645 19688
rect 172 19656 188 19658
rect 122 19640 188 19656
rect 1650 19594 1716 19610
rect 1650 19592 1666 19594
rect 193 19562 219 19592
rect 1619 19562 1666 19592
rect 122 19498 188 19514
rect 122 19464 138 19498
rect 172 19496 188 19498
rect 1650 19560 1666 19562
rect 1700 19560 1716 19594
rect 1650 19544 1716 19560
rect 172 19466 219 19496
rect 1619 19466 1645 19496
rect 172 19464 188 19466
rect 122 19448 188 19464
rect 1650 19402 1716 19418
rect 1650 19400 1666 19402
rect 193 19370 219 19400
rect 1619 19370 1666 19400
rect 122 19306 188 19322
rect 122 19272 138 19306
rect 172 19304 188 19306
rect 1650 19368 1666 19370
rect 1700 19368 1716 19402
rect 1650 19352 1716 19368
rect 172 19274 219 19304
rect 1619 19274 1645 19304
rect 172 19272 188 19274
rect 122 19256 188 19272
rect 1650 19210 1716 19226
rect 1650 19208 1666 19210
rect 193 19178 219 19208
rect 1619 19178 1666 19208
rect 122 19114 188 19130
rect 122 19080 138 19114
rect 172 19112 188 19114
rect 1650 19176 1666 19178
rect 1700 19176 1716 19210
rect 1650 19160 1716 19176
rect 172 19082 219 19112
rect 1619 19082 1645 19112
rect 172 19080 188 19082
rect 122 19064 188 19080
rect 1650 19018 1716 19034
rect 1650 19016 1666 19018
rect 193 18986 219 19016
rect 1619 18986 1666 19016
rect 122 18922 188 18938
rect 122 18888 138 18922
rect 172 18920 188 18922
rect 1650 18984 1666 18986
rect 1700 18984 1716 19018
rect 1650 18968 1716 18984
rect 172 18890 219 18920
rect 1619 18890 1645 18920
rect 172 18888 188 18890
rect 122 18872 188 18888
rect 1650 18826 1716 18842
rect 1650 18824 1666 18826
rect 193 18794 219 18824
rect 1619 18794 1666 18824
rect 122 18730 188 18746
rect 122 18696 138 18730
rect 172 18728 188 18730
rect 1650 18792 1666 18794
rect 1700 18792 1716 18826
rect 1650 18776 1716 18792
rect 172 18698 219 18728
rect 1619 18698 1645 18728
rect 172 18696 188 18698
rect 122 18680 188 18696
rect 1650 18634 1716 18650
rect 1650 18632 1666 18634
rect 193 18602 219 18632
rect 1619 18602 1666 18632
rect 122 18538 188 18554
rect 122 18504 138 18538
rect 172 18536 188 18538
rect 1650 18600 1666 18602
rect 1700 18600 1716 18634
rect 1650 18584 1716 18600
rect 172 18506 219 18536
rect 1619 18506 1645 18536
rect 172 18504 188 18506
rect 122 18488 188 18504
rect 1650 18442 1716 18458
rect 1650 18440 1666 18442
rect 193 18410 219 18440
rect 1619 18410 1666 18440
rect 122 18346 188 18362
rect 122 18312 138 18346
rect 172 18344 188 18346
rect 1650 18408 1666 18410
rect 1700 18408 1716 18442
rect 1650 18392 1716 18408
rect 172 18314 219 18344
rect 1619 18314 1645 18344
rect 172 18312 188 18314
rect 122 18296 188 18312
rect 1650 18250 1716 18266
rect 1650 18248 1666 18250
rect 193 18218 219 18248
rect 1619 18218 1666 18248
rect 122 18154 188 18170
rect 122 18120 138 18154
rect 172 18152 188 18154
rect 1650 18216 1666 18218
rect 1700 18216 1716 18250
rect 1650 18200 1716 18216
rect 172 18122 219 18152
rect 1619 18122 1645 18152
rect 172 18120 188 18122
rect 122 18104 188 18120
rect 1650 18058 1716 18074
rect 1650 18056 1666 18058
rect 193 18026 219 18056
rect 1619 18026 1666 18056
rect 122 17962 188 17978
rect 122 17928 138 17962
rect 172 17960 188 17962
rect 1650 18024 1666 18026
rect 1700 18024 1716 18058
rect 1650 18008 1716 18024
rect 172 17930 219 17960
rect 1619 17930 1645 17960
rect 172 17928 188 17930
rect 122 17912 188 17928
rect 1650 17866 1716 17882
rect 1650 17864 1666 17866
rect 193 17834 219 17864
rect 1619 17834 1666 17864
rect 122 17770 188 17786
rect 122 17736 138 17770
rect 172 17768 188 17770
rect 1650 17832 1666 17834
rect 1700 17832 1716 17866
rect 1650 17816 1716 17832
rect 172 17738 219 17768
rect 1619 17738 1645 17768
rect 172 17736 188 17738
rect 122 17720 188 17736
rect 1650 17674 1716 17690
rect 1650 17672 1666 17674
rect 193 17642 219 17672
rect 1619 17642 1666 17672
rect 122 17578 188 17594
rect 122 17544 138 17578
rect 172 17576 188 17578
rect 1650 17640 1666 17642
rect 1700 17640 1716 17674
rect 1650 17624 1716 17640
rect 172 17546 219 17576
rect 1619 17546 1645 17576
rect 172 17544 188 17546
rect 122 17528 188 17544
rect 1650 17482 1716 17498
rect 1650 17480 1666 17482
rect 193 17450 219 17480
rect 1619 17450 1666 17480
rect 122 17386 188 17402
rect 122 17352 138 17386
rect 172 17384 188 17386
rect 1650 17448 1666 17450
rect 1700 17448 1716 17482
rect 1650 17432 1716 17448
rect 172 17354 219 17384
rect 1619 17354 1645 17384
rect 172 17352 188 17354
rect 122 17336 188 17352
rect 1650 17290 1716 17306
rect 1650 17288 1666 17290
rect 193 17258 219 17288
rect 1619 17258 1666 17288
rect 122 17194 188 17210
rect 122 17160 138 17194
rect 172 17192 188 17194
rect 1650 17256 1666 17258
rect 1700 17256 1716 17290
rect 1650 17240 1716 17256
rect 172 17162 219 17192
rect 1619 17162 1645 17192
rect 172 17160 188 17162
rect 122 17144 188 17160
rect 1650 17098 1716 17114
rect 1650 17096 1666 17098
rect 193 17066 219 17096
rect 1619 17066 1666 17096
rect 122 17002 188 17018
rect 122 16968 138 17002
rect 172 17000 188 17002
rect 1650 17064 1666 17066
rect 1700 17064 1716 17098
rect 1650 17048 1716 17064
rect 172 16970 219 17000
rect 1619 16970 1645 17000
rect 172 16968 188 16970
rect 122 16952 188 16968
rect 1650 16906 1716 16922
rect 1650 16904 1666 16906
rect 193 16874 219 16904
rect 1619 16874 1666 16904
rect 122 16810 188 16826
rect 122 16776 138 16810
rect 172 16808 188 16810
rect 1650 16872 1666 16874
rect 1700 16872 1716 16906
rect 1650 16856 1716 16872
rect 172 16778 219 16808
rect 1619 16778 1645 16808
rect 172 16776 188 16778
rect 122 16760 188 16776
rect 1650 16714 1716 16730
rect 1650 16712 1666 16714
rect 193 16682 219 16712
rect 1619 16682 1666 16712
rect 122 16618 188 16634
rect 122 16584 138 16618
rect 172 16616 188 16618
rect 1650 16680 1666 16682
rect 1700 16680 1716 16714
rect 1650 16664 1716 16680
rect 172 16586 219 16616
rect 1619 16586 1645 16616
rect 172 16584 188 16586
rect 122 16568 188 16584
rect 1650 16522 1716 16538
rect 1650 16520 1666 16522
rect 193 16490 219 16520
rect 1619 16490 1666 16520
rect 122 16426 188 16442
rect 122 16392 138 16426
rect 172 16424 188 16426
rect 1650 16488 1666 16490
rect 1700 16488 1716 16522
rect 1650 16472 1716 16488
rect 172 16394 219 16424
rect 1619 16394 1645 16424
rect 172 16392 188 16394
rect 122 16376 188 16392
rect 1650 16330 1716 16346
rect 1650 16328 1666 16330
rect 193 16298 219 16328
rect 1619 16298 1666 16328
rect 122 16234 188 16250
rect 122 16200 138 16234
rect 172 16232 188 16234
rect 1650 16296 1666 16298
rect 1700 16296 1716 16330
rect 1650 16280 1716 16296
rect 172 16202 219 16232
rect 1619 16202 1645 16232
rect 172 16200 188 16202
rect 122 16184 188 16200
rect 1650 16138 1716 16154
rect 1650 16136 1666 16138
rect 193 16106 219 16136
rect 1619 16106 1666 16136
rect 122 16042 188 16058
rect 122 16008 138 16042
rect 172 16040 188 16042
rect 1650 16104 1666 16106
rect 1700 16104 1716 16138
rect 1650 16088 1716 16104
rect 172 16010 219 16040
rect 1619 16010 1645 16040
rect 172 16008 188 16010
rect 122 15992 188 16008
rect 1650 15946 1716 15962
rect 1650 15944 1666 15946
rect 193 15914 219 15944
rect 1619 15914 1666 15944
rect 122 15850 188 15866
rect 122 15816 138 15850
rect 172 15848 188 15850
rect 1650 15912 1666 15914
rect 1700 15912 1716 15946
rect 1650 15896 1716 15912
rect 172 15818 219 15848
rect 1619 15818 1645 15848
rect 172 15816 188 15818
rect 122 15800 188 15816
rect 1650 15754 1716 15770
rect 1650 15752 1666 15754
rect 193 15722 219 15752
rect 1619 15722 1666 15752
rect 122 15658 188 15674
rect 122 15624 138 15658
rect 172 15656 188 15658
rect 1650 15720 1666 15722
rect 1700 15720 1716 15754
rect 1650 15704 1716 15720
rect 172 15626 219 15656
rect 1619 15626 1645 15656
rect 172 15624 188 15626
rect 122 15608 188 15624
rect 1650 15562 1716 15578
rect 1650 15560 1666 15562
rect 193 15530 219 15560
rect 1619 15530 1666 15560
rect 122 15466 188 15482
rect 122 15432 138 15466
rect 172 15464 188 15466
rect 1650 15528 1666 15530
rect 1700 15528 1716 15562
rect 1650 15512 1716 15528
rect 172 15434 219 15464
rect 1619 15434 1645 15464
rect 172 15432 188 15434
rect 122 15416 188 15432
rect 1650 15370 1716 15386
rect 1650 15368 1666 15370
rect 193 15338 219 15368
rect 1619 15338 1666 15368
rect 122 15274 188 15290
rect 122 15240 138 15274
rect 172 15272 188 15274
rect 1650 15336 1666 15338
rect 1700 15336 1716 15370
rect 1650 15320 1716 15336
rect 172 15242 219 15272
rect 1619 15242 1645 15272
rect 172 15240 188 15242
rect 122 15224 188 15240
rect 1650 15178 1716 15194
rect 1650 15176 1666 15178
rect 193 15146 219 15176
rect 1619 15146 1666 15176
rect 122 15082 188 15098
rect 122 15048 138 15082
rect 172 15080 188 15082
rect 1650 15144 1666 15146
rect 1700 15144 1716 15178
rect 1650 15128 1716 15144
rect 172 15050 219 15080
rect 1619 15050 1645 15080
rect 172 15048 188 15050
rect 122 15032 188 15048
rect 1650 14986 1716 15002
rect 1650 14984 1666 14986
rect 193 14954 219 14984
rect 1619 14954 1666 14984
rect 122 14890 188 14906
rect 122 14856 138 14890
rect 172 14888 188 14890
rect 1650 14952 1666 14954
rect 1700 14952 1716 14986
rect 1650 14936 1716 14952
rect 172 14858 219 14888
rect 1619 14858 1645 14888
rect 172 14856 188 14858
rect 122 14840 188 14856
rect 1650 14794 1716 14810
rect 1650 14792 1666 14794
rect 193 14762 219 14792
rect 1619 14762 1666 14792
rect 122 14698 188 14714
rect 122 14664 138 14698
rect 172 14696 188 14698
rect 1650 14760 1666 14762
rect 1700 14760 1716 14794
rect 1650 14744 1716 14760
rect 172 14666 219 14696
rect 1619 14666 1645 14696
rect 172 14664 188 14666
rect 122 14648 188 14664
rect 1650 14602 1716 14618
rect 1650 14600 1666 14602
rect 193 14570 219 14600
rect 1619 14570 1666 14600
rect 122 14506 188 14522
rect 122 14472 138 14506
rect 172 14504 188 14506
rect 1650 14568 1666 14570
rect 1700 14568 1716 14602
rect 1650 14552 1716 14568
rect 172 14474 219 14504
rect 1619 14474 1645 14504
rect 172 14472 188 14474
rect 122 14456 188 14472
rect 1650 14410 1716 14426
rect 1650 14408 1666 14410
rect 193 14378 219 14408
rect 1619 14378 1666 14408
rect 122 14314 188 14330
rect 122 14280 138 14314
rect 172 14312 188 14314
rect 1650 14376 1666 14378
rect 1700 14376 1716 14410
rect 1650 14360 1716 14376
rect 172 14282 219 14312
rect 1619 14282 1645 14312
rect 172 14280 188 14282
rect 122 14264 188 14280
rect 1650 14218 1716 14234
rect 1650 14216 1666 14218
rect 193 14186 219 14216
rect 1619 14186 1666 14216
rect 122 14122 188 14138
rect 122 14088 138 14122
rect 172 14120 188 14122
rect 1650 14184 1666 14186
rect 1700 14184 1716 14218
rect 1650 14168 1716 14184
rect 172 14090 219 14120
rect 1619 14090 1645 14120
rect 172 14088 188 14090
rect 122 14072 188 14088
rect 1650 14026 1716 14042
rect 1650 14024 1666 14026
rect 193 13994 219 14024
rect 1619 13994 1666 14024
rect 122 13930 188 13946
rect 122 13896 138 13930
rect 172 13928 188 13930
rect 1650 13992 1666 13994
rect 1700 13992 1716 14026
rect 1650 13976 1716 13992
rect 172 13898 219 13928
rect 1619 13898 1645 13928
rect 172 13896 188 13898
rect 122 13880 188 13896
rect 1650 13834 1716 13850
rect 1650 13832 1666 13834
rect 193 13802 219 13832
rect 1619 13802 1666 13832
rect 122 13738 188 13754
rect 122 13704 138 13738
rect 172 13736 188 13738
rect 1650 13800 1666 13802
rect 1700 13800 1716 13834
rect 1650 13784 1716 13800
rect 172 13706 219 13736
rect 1619 13706 1645 13736
rect 172 13704 188 13706
rect 122 13688 188 13704
rect 1650 13642 1716 13658
rect 1650 13640 1666 13642
rect 193 13610 219 13640
rect 1619 13610 1666 13640
rect 122 13546 188 13562
rect 122 13512 138 13546
rect 172 13544 188 13546
rect 1650 13608 1666 13610
rect 1700 13608 1716 13642
rect 1650 13592 1716 13608
rect 172 13514 219 13544
rect 1619 13514 1645 13544
rect 172 13512 188 13514
rect 122 13496 188 13512
rect 1650 13450 1716 13466
rect 1650 13448 1666 13450
rect 193 13418 219 13448
rect 1619 13418 1666 13448
rect 122 13354 188 13370
rect 122 13320 138 13354
rect 172 13352 188 13354
rect 1650 13416 1666 13418
rect 1700 13416 1716 13450
rect 1650 13400 1716 13416
rect 172 13322 219 13352
rect 1619 13322 1645 13352
rect 172 13320 188 13322
rect 122 13304 188 13320
rect 1650 13258 1716 13274
rect 1650 13256 1666 13258
rect 193 13226 219 13256
rect 1619 13226 1666 13256
rect 122 13162 188 13178
rect 122 13128 138 13162
rect 172 13160 188 13162
rect 1650 13224 1666 13226
rect 1700 13224 1716 13258
rect 1650 13208 1716 13224
rect 172 13130 219 13160
rect 1619 13130 1645 13160
rect 172 13128 188 13130
rect 122 13112 188 13128
rect 1650 13066 1716 13082
rect 1650 13064 1666 13066
rect 193 13034 219 13064
rect 1619 13034 1666 13064
rect 122 12970 188 12986
rect 122 12936 138 12970
rect 172 12968 188 12970
rect 1650 13032 1666 13034
rect 1700 13032 1716 13066
rect 1650 13016 1716 13032
rect 172 12938 219 12968
rect 1619 12938 1645 12968
rect 172 12936 188 12938
rect 122 12920 188 12936
rect 1650 12874 1716 12890
rect 1650 12872 1666 12874
rect 193 12842 219 12872
rect 1619 12842 1666 12872
rect 122 12778 188 12794
rect 122 12744 138 12778
rect 172 12776 188 12778
rect 1650 12840 1666 12842
rect 1700 12840 1716 12874
rect 1650 12824 1716 12840
rect 172 12746 219 12776
rect 1619 12746 1645 12776
rect 172 12744 188 12746
rect 122 12728 188 12744
rect 1650 12682 1716 12698
rect 1650 12680 1666 12682
rect 193 12650 219 12680
rect 1619 12650 1666 12680
rect 122 12586 188 12602
rect 122 12552 138 12586
rect 172 12584 188 12586
rect 1650 12648 1666 12650
rect 1700 12648 1716 12682
rect 1650 12632 1716 12648
rect 172 12554 219 12584
rect 1619 12554 1645 12584
rect 172 12552 188 12554
rect 122 12536 188 12552
rect 1650 12490 1716 12506
rect 1650 12488 1666 12490
rect 193 12458 219 12488
rect 1619 12458 1666 12488
rect 122 12394 188 12410
rect 122 12360 138 12394
rect 172 12392 188 12394
rect 1650 12456 1666 12458
rect 1700 12456 1716 12490
rect 1650 12440 1716 12456
rect 172 12362 219 12392
rect 1619 12362 1645 12392
rect 172 12360 188 12362
rect 122 12344 188 12360
rect 1650 12298 1716 12314
rect 1650 12296 1666 12298
rect 193 12266 219 12296
rect 1619 12266 1666 12296
rect 122 12202 188 12218
rect 122 12168 138 12202
rect 172 12200 188 12202
rect 1650 12264 1666 12266
rect 1700 12264 1716 12298
rect 1650 12248 1716 12264
rect 172 12170 219 12200
rect 1619 12170 1645 12200
rect 172 12168 188 12170
rect 122 12152 188 12168
rect 1650 12106 1716 12122
rect 1650 12104 1666 12106
rect 193 12074 219 12104
rect 1619 12074 1666 12104
rect 122 12010 188 12026
rect 122 11976 138 12010
rect 172 12008 188 12010
rect 1650 12072 1666 12074
rect 1700 12072 1716 12106
rect 1650 12056 1716 12072
rect 172 11978 219 12008
rect 1619 11978 1645 12008
rect 172 11976 188 11978
rect 122 11960 188 11976
rect 1650 11914 1716 11930
rect 1650 11912 1666 11914
rect 193 11882 219 11912
rect 1619 11882 1666 11912
rect 122 11818 188 11834
rect 122 11784 138 11818
rect 172 11816 188 11818
rect 1650 11880 1666 11882
rect 1700 11880 1716 11914
rect 1650 11864 1716 11880
rect 172 11786 219 11816
rect 1619 11786 1645 11816
rect 172 11784 188 11786
rect 122 11768 188 11784
rect 1650 11722 1716 11738
rect 1650 11720 1666 11722
rect 193 11690 219 11720
rect 1619 11690 1666 11720
rect 122 11626 188 11642
rect 122 11592 138 11626
rect 172 11624 188 11626
rect 1650 11688 1666 11690
rect 1700 11688 1716 11722
rect 1650 11672 1716 11688
rect 172 11594 219 11624
rect 1619 11594 1645 11624
rect 172 11592 188 11594
rect 122 11576 188 11592
rect 1650 11530 1716 11546
rect 1650 11528 1666 11530
rect 193 11498 219 11528
rect 1619 11498 1666 11528
rect 122 11434 188 11450
rect 122 11400 138 11434
rect 172 11432 188 11434
rect 1650 11496 1666 11498
rect 1700 11496 1716 11530
rect 1650 11480 1716 11496
rect 172 11402 219 11432
rect 1619 11402 1645 11432
rect 172 11400 188 11402
rect 122 11384 188 11400
rect 1650 11338 1716 11354
rect 1650 11336 1666 11338
rect 193 11306 219 11336
rect 1619 11306 1666 11336
rect 122 11242 188 11258
rect 122 11208 138 11242
rect 172 11240 188 11242
rect 1650 11304 1666 11306
rect 1700 11304 1716 11338
rect 1650 11288 1716 11304
rect 172 11210 219 11240
rect 1619 11210 1645 11240
rect 172 11208 188 11210
rect 122 11192 188 11208
rect 1650 11146 1716 11162
rect 1650 11144 1666 11146
rect 193 11114 219 11144
rect 1619 11114 1666 11144
rect 122 11050 188 11066
rect 122 11016 138 11050
rect 172 11048 188 11050
rect 1650 11112 1666 11114
rect 1700 11112 1716 11146
rect 1650 11096 1716 11112
rect 172 11018 219 11048
rect 1619 11018 1645 11048
rect 172 11016 188 11018
rect 122 11000 188 11016
rect 1650 10954 1716 10970
rect 1650 10952 1666 10954
rect 193 10922 219 10952
rect 1619 10922 1666 10952
rect 122 10858 188 10874
rect 122 10824 138 10858
rect 172 10856 188 10858
rect 1650 10920 1666 10922
rect 1700 10920 1716 10954
rect 1650 10904 1716 10920
rect 172 10826 219 10856
rect 1619 10826 1645 10856
rect 172 10824 188 10826
rect 122 10808 188 10824
rect 1650 10762 1716 10778
rect 1650 10760 1666 10762
rect 193 10730 219 10760
rect 1619 10730 1666 10760
rect 122 10666 188 10682
rect 122 10632 138 10666
rect 172 10664 188 10666
rect 1650 10728 1666 10730
rect 1700 10728 1716 10762
rect 1650 10712 1716 10728
rect 172 10634 219 10664
rect 1619 10634 1645 10664
rect 172 10632 188 10634
rect 122 10616 188 10632
rect 1650 10570 1716 10586
rect 1650 10568 1666 10570
rect 193 10538 219 10568
rect 1619 10538 1666 10568
rect 122 10474 188 10490
rect 122 10440 138 10474
rect 172 10472 188 10474
rect 1650 10536 1666 10538
rect 1700 10536 1716 10570
rect 1650 10520 1716 10536
rect 172 10442 219 10472
rect 1619 10442 1645 10472
rect 172 10440 188 10442
rect 122 10424 188 10440
rect 1650 10378 1716 10394
rect 1650 10376 1666 10378
rect 193 10346 219 10376
rect 1619 10346 1666 10376
rect 122 10282 188 10298
rect 122 10248 138 10282
rect 172 10280 188 10282
rect 1650 10344 1666 10346
rect 1700 10344 1716 10378
rect 1650 10328 1716 10344
rect 172 10250 219 10280
rect 1619 10250 1645 10280
rect 172 10248 188 10250
rect 122 10232 188 10248
rect 1650 10186 1716 10202
rect 1650 10184 1666 10186
rect 193 10154 219 10184
rect 1619 10154 1666 10184
rect 122 10090 188 10106
rect 122 10056 138 10090
rect 172 10088 188 10090
rect 1650 10152 1666 10154
rect 1700 10152 1716 10186
rect 1650 10136 1716 10152
rect 172 10058 219 10088
rect 1619 10058 1645 10088
rect 172 10056 188 10058
rect 122 10040 188 10056
rect 1650 9994 1716 10010
rect 1650 9992 1666 9994
rect 193 9962 219 9992
rect 1619 9962 1666 9992
rect 122 9898 188 9914
rect 122 9864 138 9898
rect 172 9896 188 9898
rect 1650 9960 1666 9962
rect 1700 9960 1716 9994
rect 1650 9944 1716 9960
rect 172 9866 219 9896
rect 1619 9866 1645 9896
rect 172 9864 188 9866
rect 122 9848 188 9864
rect 1650 9802 1716 9818
rect 1650 9800 1666 9802
rect 193 9770 219 9800
rect 1619 9770 1666 9800
rect 122 9706 188 9722
rect 122 9672 138 9706
rect 172 9704 188 9706
rect 1650 9768 1666 9770
rect 1700 9768 1716 9802
rect 1650 9752 1716 9768
rect 172 9674 219 9704
rect 1619 9674 1645 9704
rect 172 9672 188 9674
rect 122 9656 188 9672
rect 1650 9610 1716 9626
rect 1650 9608 1666 9610
rect 193 9578 219 9608
rect 1619 9578 1666 9608
rect 122 9514 188 9530
rect 122 9480 138 9514
rect 172 9512 188 9514
rect 1650 9576 1666 9578
rect 1700 9576 1716 9610
rect 1650 9560 1716 9576
rect 172 9482 219 9512
rect 1619 9482 1645 9512
rect 172 9480 188 9482
rect 122 9464 188 9480
rect 1650 9418 1716 9434
rect 1650 9416 1666 9418
rect 193 9386 219 9416
rect 1619 9386 1666 9416
rect 122 9322 188 9338
rect 122 9288 138 9322
rect 172 9320 188 9322
rect 1650 9384 1666 9386
rect 1700 9384 1716 9418
rect 1650 9368 1716 9384
rect 172 9290 219 9320
rect 1619 9290 1645 9320
rect 172 9288 188 9290
rect 122 9272 188 9288
rect 1650 9226 1716 9242
rect 1650 9224 1666 9226
rect 193 9194 219 9224
rect 1619 9194 1666 9224
rect 122 9130 188 9146
rect 122 9096 138 9130
rect 172 9128 188 9130
rect 1650 9192 1666 9194
rect 1700 9192 1716 9226
rect 1650 9176 1716 9192
rect 172 9098 219 9128
rect 1619 9098 1645 9128
rect 172 9096 188 9098
rect 122 9080 188 9096
rect 1650 9034 1716 9050
rect 1650 9032 1666 9034
rect 193 9002 219 9032
rect 1619 9002 1666 9032
rect 122 8938 188 8954
rect 122 8904 138 8938
rect 172 8936 188 8938
rect 1650 9000 1666 9002
rect 1700 9000 1716 9034
rect 1650 8984 1716 9000
rect 172 8906 219 8936
rect 1619 8906 1645 8936
rect 172 8904 188 8906
rect 122 8888 188 8904
rect 1650 8842 1716 8858
rect 1650 8840 1666 8842
rect 193 8810 219 8840
rect 1619 8810 1666 8840
rect 122 8746 188 8762
rect 122 8712 138 8746
rect 172 8744 188 8746
rect 1650 8808 1666 8810
rect 1700 8808 1716 8842
rect 1650 8792 1716 8808
rect 172 8714 219 8744
rect 1619 8714 1645 8744
rect 172 8712 188 8714
rect 122 8696 188 8712
rect 1650 8650 1716 8666
rect 1650 8648 1666 8650
rect 193 8618 219 8648
rect 1619 8618 1666 8648
rect 122 8554 188 8570
rect 122 8520 138 8554
rect 172 8552 188 8554
rect 1650 8616 1666 8618
rect 1700 8616 1716 8650
rect 1650 8600 1716 8616
rect 172 8522 219 8552
rect 1619 8522 1645 8552
rect 172 8520 188 8522
rect 122 8504 188 8520
rect 1650 8458 1716 8474
rect 1650 8456 1666 8458
rect 193 8426 219 8456
rect 1619 8426 1666 8456
rect 122 8362 188 8378
rect 122 8328 138 8362
rect 172 8360 188 8362
rect 1650 8424 1666 8426
rect 1700 8424 1716 8458
rect 1650 8408 1716 8424
rect 172 8330 219 8360
rect 1619 8330 1645 8360
rect 172 8328 188 8330
rect 122 8312 188 8328
rect 1650 8266 1716 8282
rect 1650 8264 1666 8266
rect 193 8234 219 8264
rect 1619 8234 1666 8264
rect 122 8170 188 8186
rect 122 8136 138 8170
rect 172 8168 188 8170
rect 1650 8232 1666 8234
rect 1700 8232 1716 8266
rect 1650 8216 1716 8232
rect 172 8138 219 8168
rect 1619 8138 1645 8168
rect 172 8136 188 8138
rect 122 8120 188 8136
rect 1650 8074 1716 8090
rect 1650 8072 1666 8074
rect 193 8042 219 8072
rect 1619 8042 1666 8072
rect 122 7978 188 7994
rect 122 7944 138 7978
rect 172 7976 188 7978
rect 1650 8040 1666 8042
rect 1700 8040 1716 8074
rect 1650 8024 1716 8040
rect 172 7946 219 7976
rect 1619 7946 1645 7976
rect 172 7944 188 7946
rect 122 7928 188 7944
rect 1650 7882 1716 7898
rect 1650 7880 1666 7882
rect 193 7850 219 7880
rect 1619 7850 1666 7880
rect 122 7786 188 7802
rect 122 7752 138 7786
rect 172 7784 188 7786
rect 1650 7848 1666 7850
rect 1700 7848 1716 7882
rect 1650 7832 1716 7848
rect 172 7754 219 7784
rect 1619 7754 1645 7784
rect 172 7752 188 7754
rect 122 7736 188 7752
rect 1650 7690 1716 7706
rect 1650 7688 1666 7690
rect 193 7658 219 7688
rect 1619 7658 1666 7688
rect 122 7594 188 7610
rect 122 7560 138 7594
rect 172 7592 188 7594
rect 1650 7656 1666 7658
rect 1700 7656 1716 7690
rect 1650 7640 1716 7656
rect 172 7562 219 7592
rect 1619 7562 1645 7592
rect 172 7560 188 7562
rect 122 7544 188 7560
rect 1650 7498 1716 7514
rect 1650 7496 1666 7498
rect 193 7466 219 7496
rect 1619 7466 1666 7496
rect 122 7402 188 7418
rect 122 7368 138 7402
rect 172 7400 188 7402
rect 1650 7464 1666 7466
rect 1700 7464 1716 7498
rect 1650 7448 1716 7464
rect 172 7370 219 7400
rect 1619 7370 1645 7400
rect 172 7368 188 7370
rect 122 7352 188 7368
rect 1650 7306 1716 7322
rect 1650 7304 1666 7306
rect 193 7274 219 7304
rect 1619 7274 1666 7304
rect 122 7210 188 7226
rect 122 7176 138 7210
rect 172 7208 188 7210
rect 1650 7272 1666 7274
rect 1700 7272 1716 7306
rect 1650 7256 1716 7272
rect 172 7178 219 7208
rect 1619 7178 1645 7208
rect 172 7176 188 7178
rect 122 7160 188 7176
rect 1650 7114 1716 7130
rect 1650 7112 1666 7114
rect 193 7082 219 7112
rect 1619 7082 1666 7112
rect 122 7018 188 7034
rect 122 6984 138 7018
rect 172 7016 188 7018
rect 1650 7080 1666 7082
rect 1700 7080 1716 7114
rect 1650 7064 1716 7080
rect 172 6986 219 7016
rect 1619 6986 1645 7016
rect 172 6984 188 6986
rect 122 6968 188 6984
rect 1650 6922 1716 6938
rect 1650 6920 1666 6922
rect 193 6890 219 6920
rect 1619 6890 1666 6920
rect 122 6826 188 6842
rect 122 6792 138 6826
rect 172 6824 188 6826
rect 1650 6888 1666 6890
rect 1700 6888 1716 6922
rect 1650 6872 1716 6888
rect 172 6794 219 6824
rect 1619 6794 1645 6824
rect 172 6792 188 6794
rect 122 6776 188 6792
rect 1650 6730 1716 6746
rect 1650 6728 1666 6730
rect 193 6698 219 6728
rect 1619 6698 1666 6728
rect 122 6634 188 6650
rect 122 6600 138 6634
rect 172 6632 188 6634
rect 1650 6696 1666 6698
rect 1700 6696 1716 6730
rect 1650 6680 1716 6696
rect 172 6602 219 6632
rect 1619 6602 1645 6632
rect 172 6600 188 6602
rect 122 6584 188 6600
rect 1650 6538 1716 6554
rect 1650 6536 1666 6538
rect 193 6506 219 6536
rect 1619 6506 1666 6536
rect 122 6442 188 6458
rect 122 6408 138 6442
rect 172 6440 188 6442
rect 1650 6504 1666 6506
rect 1700 6504 1716 6538
rect 1650 6488 1716 6504
rect 172 6410 219 6440
rect 1619 6410 1645 6440
rect 172 6408 188 6410
rect 122 6392 188 6408
rect 1650 6346 1716 6362
rect 1650 6344 1666 6346
rect 193 6314 219 6344
rect 1619 6314 1666 6344
rect 122 6250 188 6266
rect 122 6216 138 6250
rect 172 6248 188 6250
rect 1650 6312 1666 6314
rect 1700 6312 1716 6346
rect 1650 6296 1716 6312
rect 172 6218 219 6248
rect 1619 6218 1645 6248
rect 172 6216 188 6218
rect 122 6200 188 6216
rect 1650 6154 1716 6170
rect 1650 6152 1666 6154
rect 193 6122 219 6152
rect 1619 6122 1666 6152
rect 122 6058 188 6074
rect 122 6024 138 6058
rect 172 6056 188 6058
rect 1650 6120 1666 6122
rect 1700 6120 1716 6154
rect 1650 6104 1716 6120
rect 172 6026 219 6056
rect 1619 6026 1645 6056
rect 172 6024 188 6026
rect 122 6008 188 6024
rect 1650 5962 1716 5978
rect 1650 5960 1666 5962
rect 193 5930 219 5960
rect 1619 5930 1666 5960
rect 122 5866 188 5882
rect 122 5832 138 5866
rect 172 5864 188 5866
rect 1650 5928 1666 5930
rect 1700 5928 1716 5962
rect 1650 5912 1716 5928
rect 172 5834 219 5864
rect 1619 5834 1645 5864
rect 172 5832 188 5834
rect 122 5816 188 5832
rect 1650 5770 1716 5786
rect 1650 5768 1666 5770
rect 193 5738 219 5768
rect 1619 5738 1666 5768
rect 122 5674 188 5690
rect 122 5640 138 5674
rect 172 5672 188 5674
rect 1650 5736 1666 5738
rect 1700 5736 1716 5770
rect 1650 5720 1716 5736
rect 172 5642 219 5672
rect 1619 5642 1645 5672
rect 172 5640 188 5642
rect 122 5624 188 5640
rect 1650 5578 1716 5594
rect 1650 5576 1666 5578
rect 193 5546 219 5576
rect 1619 5546 1666 5576
rect 122 5482 188 5498
rect 122 5448 138 5482
rect 172 5480 188 5482
rect 1650 5544 1666 5546
rect 1700 5544 1716 5578
rect 1650 5528 1716 5544
rect 172 5450 219 5480
rect 1619 5450 1645 5480
rect 172 5448 188 5450
rect 122 5432 188 5448
rect 1650 5386 1716 5402
rect 1650 5384 1666 5386
rect 193 5354 219 5384
rect 1619 5354 1666 5384
rect 122 5290 188 5306
rect 122 5256 138 5290
rect 172 5288 188 5290
rect 1650 5352 1666 5354
rect 1700 5352 1716 5386
rect 1650 5336 1716 5352
rect 172 5258 219 5288
rect 1619 5258 1645 5288
rect 172 5256 188 5258
rect 122 5240 188 5256
rect 1650 5194 1716 5210
rect 1650 5192 1666 5194
rect 193 5162 219 5192
rect 1619 5162 1666 5192
rect 122 5098 188 5114
rect 122 5064 138 5098
rect 172 5096 188 5098
rect 1650 5160 1666 5162
rect 1700 5160 1716 5194
rect 1650 5144 1716 5160
rect 172 5066 219 5096
rect 1619 5066 1645 5096
rect 172 5064 188 5066
rect 122 5048 188 5064
rect 1650 5002 1716 5018
rect 1650 5000 1666 5002
rect 193 4970 219 5000
rect 1619 4970 1666 5000
rect 122 4906 188 4922
rect 122 4872 138 4906
rect 172 4904 188 4906
rect 1650 4968 1666 4970
rect 1700 4968 1716 5002
rect 1650 4952 1716 4968
rect 172 4874 219 4904
rect 1619 4874 1645 4904
rect 172 4872 188 4874
rect 122 4856 188 4872
rect 1650 4810 1716 4826
rect 1650 4808 1666 4810
rect 193 4778 219 4808
rect 1619 4778 1666 4808
rect 122 4714 188 4730
rect 122 4680 138 4714
rect 172 4712 188 4714
rect 1650 4776 1666 4778
rect 1700 4776 1716 4810
rect 1650 4760 1716 4776
rect 172 4682 219 4712
rect 1619 4682 1645 4712
rect 172 4680 188 4682
rect 122 4664 188 4680
rect 1650 4618 1716 4634
rect 1650 4616 1666 4618
rect 193 4586 219 4616
rect 1619 4586 1666 4616
rect 122 4522 188 4538
rect 122 4488 138 4522
rect 172 4520 188 4522
rect 1650 4584 1666 4586
rect 1700 4584 1716 4618
rect 1650 4568 1716 4584
rect 172 4490 219 4520
rect 1619 4490 1645 4520
rect 172 4488 188 4490
rect 122 4472 188 4488
rect 1650 4426 1716 4442
rect 1650 4424 1666 4426
rect 193 4394 219 4424
rect 1619 4394 1666 4424
rect 122 4330 188 4346
rect 122 4296 138 4330
rect 172 4328 188 4330
rect 1650 4392 1666 4394
rect 1700 4392 1716 4426
rect 1650 4376 1716 4392
rect 172 4298 219 4328
rect 1619 4298 1645 4328
rect 172 4296 188 4298
rect 122 4280 188 4296
rect 1650 4234 1716 4250
rect 1650 4232 1666 4234
rect 193 4202 219 4232
rect 1619 4202 1666 4232
rect 122 4138 188 4154
rect 122 4104 138 4138
rect 172 4136 188 4138
rect 1650 4200 1666 4202
rect 1700 4200 1716 4234
rect 1650 4184 1716 4200
rect 172 4106 219 4136
rect 1619 4106 1645 4136
rect 172 4104 188 4106
rect 122 4088 188 4104
rect 1650 4042 1716 4058
rect 1650 4040 1666 4042
rect 193 4010 219 4040
rect 1619 4010 1666 4040
rect 122 3946 188 3962
rect 122 3912 138 3946
rect 172 3944 188 3946
rect 1650 4008 1666 4010
rect 1700 4008 1716 4042
rect 1650 3992 1716 4008
rect 172 3914 219 3944
rect 1619 3914 1645 3944
rect 172 3912 188 3914
rect 122 3896 188 3912
rect 1650 3850 1716 3866
rect 1650 3848 1666 3850
rect 193 3818 219 3848
rect 1619 3818 1666 3848
rect 122 3754 188 3770
rect 122 3720 138 3754
rect 172 3752 188 3754
rect 1650 3816 1666 3818
rect 1700 3816 1716 3850
rect 1650 3800 1716 3816
rect 172 3722 219 3752
rect 1619 3722 1645 3752
rect 172 3720 188 3722
rect 122 3704 188 3720
rect 1650 3658 1716 3674
rect 1650 3656 1666 3658
rect 193 3626 219 3656
rect 1619 3626 1666 3656
rect 122 3562 188 3578
rect 122 3528 138 3562
rect 172 3560 188 3562
rect 1650 3624 1666 3626
rect 1700 3624 1716 3658
rect 1650 3608 1716 3624
rect 172 3530 219 3560
rect 1619 3530 1645 3560
rect 172 3528 188 3530
rect 122 3512 188 3528
rect 1650 3466 1716 3482
rect 1650 3464 1666 3466
rect 193 3434 219 3464
rect 1619 3434 1666 3464
rect 122 3370 188 3386
rect 122 3336 138 3370
rect 172 3368 188 3370
rect 1650 3432 1666 3434
rect 1700 3432 1716 3466
rect 1650 3416 1716 3432
rect 172 3338 219 3368
rect 1619 3338 1645 3368
rect 172 3336 188 3338
rect 122 3320 188 3336
rect 1650 3274 1716 3290
rect 1650 3272 1666 3274
rect 193 3242 219 3272
rect 1619 3242 1666 3272
rect 122 3178 188 3194
rect 122 3144 138 3178
rect 172 3176 188 3178
rect 1650 3240 1666 3242
rect 1700 3240 1716 3274
rect 1650 3224 1716 3240
rect 172 3146 219 3176
rect 1619 3146 1645 3176
rect 172 3144 188 3146
rect 122 3128 188 3144
rect 1650 3082 1716 3098
rect 1650 3080 1666 3082
rect 193 3050 219 3080
rect 1619 3050 1666 3080
rect 122 2986 188 3002
rect 122 2952 138 2986
rect 172 2984 188 2986
rect 1650 3048 1666 3050
rect 1700 3048 1716 3082
rect 1650 3032 1716 3048
rect 172 2954 219 2984
rect 1619 2954 1645 2984
rect 172 2952 188 2954
rect 122 2936 188 2952
rect 1650 2890 1716 2906
rect 1650 2888 1666 2890
rect 193 2858 219 2888
rect 1619 2858 1666 2888
rect 122 2794 188 2810
rect 122 2760 138 2794
rect 172 2792 188 2794
rect 1650 2856 1666 2858
rect 1700 2856 1716 2890
rect 1650 2840 1716 2856
rect 172 2762 219 2792
rect 1619 2762 1645 2792
rect 172 2760 188 2762
rect 122 2744 188 2760
rect 1650 2698 1716 2714
rect 1650 2696 1666 2698
rect 193 2666 219 2696
rect 1619 2666 1666 2696
rect 122 2602 188 2618
rect 122 2568 138 2602
rect 172 2600 188 2602
rect 1650 2664 1666 2666
rect 1700 2664 1716 2698
rect 1650 2648 1716 2664
rect 172 2570 219 2600
rect 1619 2570 1645 2600
rect 172 2568 188 2570
rect 122 2552 188 2568
rect 1650 2506 1716 2522
rect 1650 2504 1666 2506
rect 193 2474 219 2504
rect 1619 2474 1666 2504
rect 122 2410 188 2426
rect 122 2376 138 2410
rect 172 2408 188 2410
rect 1650 2472 1666 2474
rect 1700 2472 1716 2506
rect 1650 2456 1716 2472
rect 172 2378 219 2408
rect 1619 2378 1645 2408
rect 172 2376 188 2378
rect 122 2360 188 2376
rect 1650 2314 1716 2330
rect 1650 2312 1666 2314
rect 193 2282 219 2312
rect 1619 2282 1666 2312
rect 122 2218 188 2234
rect 122 2184 138 2218
rect 172 2216 188 2218
rect 1650 2280 1666 2282
rect 1700 2280 1716 2314
rect 1650 2264 1716 2280
rect 172 2186 219 2216
rect 1619 2186 1645 2216
rect 172 2184 188 2186
rect 122 2168 188 2184
rect 1650 2122 1716 2138
rect 1650 2120 1666 2122
rect 193 2090 219 2120
rect 1619 2090 1666 2120
rect 122 2026 188 2042
rect 122 1992 138 2026
rect 172 2024 188 2026
rect 1650 2088 1666 2090
rect 1700 2088 1716 2122
rect 1650 2072 1716 2088
rect 172 1994 219 2024
rect 1619 1994 1645 2024
rect 172 1992 188 1994
rect 122 1976 188 1992
rect 1650 1930 1716 1946
rect 1650 1928 1666 1930
rect 193 1898 219 1928
rect 1619 1898 1666 1928
rect 122 1834 188 1850
rect 122 1800 138 1834
rect 172 1832 188 1834
rect 1650 1896 1666 1898
rect 1700 1896 1716 1930
rect 1650 1880 1716 1896
rect 172 1802 219 1832
rect 1619 1802 1645 1832
rect 172 1800 188 1802
rect 122 1784 188 1800
rect 1650 1738 1716 1754
rect 1650 1736 1666 1738
rect 193 1706 219 1736
rect 1619 1706 1666 1736
rect 122 1642 188 1658
rect 122 1608 138 1642
rect 172 1640 188 1642
rect 1650 1704 1666 1706
rect 1700 1704 1716 1738
rect 1650 1688 1716 1704
rect 172 1610 219 1640
rect 1619 1610 1645 1640
rect 172 1608 188 1610
rect 122 1592 188 1608
rect 1650 1546 1716 1562
rect 1650 1544 1666 1546
rect 193 1514 219 1544
rect 1619 1514 1666 1544
rect 122 1450 188 1466
rect 122 1416 138 1450
rect 172 1448 188 1450
rect 1650 1512 1666 1514
rect 1700 1512 1716 1546
rect 1650 1496 1716 1512
rect 172 1418 219 1448
rect 1619 1418 1645 1448
rect 172 1416 188 1418
rect 122 1400 188 1416
rect 1650 1354 1716 1370
rect 1650 1352 1666 1354
rect 193 1322 219 1352
rect 1619 1322 1666 1352
rect 122 1258 188 1274
rect 122 1224 138 1258
rect 172 1256 188 1258
rect 1650 1320 1666 1322
rect 1700 1320 1716 1354
rect 1650 1304 1716 1320
rect 172 1226 219 1256
rect 1619 1226 1645 1256
rect 172 1224 188 1226
rect 122 1208 188 1224
rect 1650 1162 1716 1178
rect 1650 1160 1666 1162
rect 193 1130 219 1160
rect 1619 1130 1666 1160
rect 122 1066 188 1082
rect 122 1032 138 1066
rect 172 1064 188 1066
rect 1650 1128 1666 1130
rect 1700 1128 1716 1162
rect 1650 1112 1716 1128
rect 172 1034 219 1064
rect 1619 1034 1645 1064
rect 172 1032 188 1034
rect 122 1016 188 1032
rect 1650 970 1716 986
rect 1650 968 1666 970
rect 193 938 219 968
rect 1619 938 1666 968
rect 122 874 188 890
rect 122 840 138 874
rect 172 872 188 874
rect 1650 936 1666 938
rect 1700 936 1716 970
rect 1650 920 1716 936
rect 172 842 219 872
rect 1619 842 1645 872
rect 172 840 188 842
rect 122 824 188 840
rect 1650 778 1716 794
rect 1650 776 1666 778
rect 193 746 219 776
rect 1619 746 1666 776
rect 1650 744 1666 746
rect 1700 744 1716 778
rect 1650 728 1716 744
<< polycont >>
rect 138 21768 172 21802
rect 138 21576 172 21610
rect 1666 21672 1700 21706
rect 138 21384 172 21418
rect 1666 21480 1700 21514
rect 138 21192 172 21226
rect 1666 21288 1700 21322
rect 138 21000 172 21034
rect 1666 21096 1700 21130
rect 138 20808 172 20842
rect 1666 20904 1700 20938
rect 138 20616 172 20650
rect 1666 20712 1700 20746
rect 138 20424 172 20458
rect 1666 20520 1700 20554
rect 138 20232 172 20266
rect 1666 20328 1700 20362
rect 138 20040 172 20074
rect 1666 20136 1700 20170
rect 138 19848 172 19882
rect 1666 19944 1700 19978
rect 138 19656 172 19690
rect 1666 19752 1700 19786
rect 138 19464 172 19498
rect 1666 19560 1700 19594
rect 138 19272 172 19306
rect 1666 19368 1700 19402
rect 138 19080 172 19114
rect 1666 19176 1700 19210
rect 138 18888 172 18922
rect 1666 18984 1700 19018
rect 138 18696 172 18730
rect 1666 18792 1700 18826
rect 138 18504 172 18538
rect 1666 18600 1700 18634
rect 138 18312 172 18346
rect 1666 18408 1700 18442
rect 138 18120 172 18154
rect 1666 18216 1700 18250
rect 138 17928 172 17962
rect 1666 18024 1700 18058
rect 138 17736 172 17770
rect 1666 17832 1700 17866
rect 138 17544 172 17578
rect 1666 17640 1700 17674
rect 138 17352 172 17386
rect 1666 17448 1700 17482
rect 138 17160 172 17194
rect 1666 17256 1700 17290
rect 138 16968 172 17002
rect 1666 17064 1700 17098
rect 138 16776 172 16810
rect 1666 16872 1700 16906
rect 138 16584 172 16618
rect 1666 16680 1700 16714
rect 138 16392 172 16426
rect 1666 16488 1700 16522
rect 138 16200 172 16234
rect 1666 16296 1700 16330
rect 138 16008 172 16042
rect 1666 16104 1700 16138
rect 138 15816 172 15850
rect 1666 15912 1700 15946
rect 138 15624 172 15658
rect 1666 15720 1700 15754
rect 138 15432 172 15466
rect 1666 15528 1700 15562
rect 138 15240 172 15274
rect 1666 15336 1700 15370
rect 138 15048 172 15082
rect 1666 15144 1700 15178
rect 138 14856 172 14890
rect 1666 14952 1700 14986
rect 138 14664 172 14698
rect 1666 14760 1700 14794
rect 138 14472 172 14506
rect 1666 14568 1700 14602
rect 138 14280 172 14314
rect 1666 14376 1700 14410
rect 138 14088 172 14122
rect 1666 14184 1700 14218
rect 138 13896 172 13930
rect 1666 13992 1700 14026
rect 138 13704 172 13738
rect 1666 13800 1700 13834
rect 138 13512 172 13546
rect 1666 13608 1700 13642
rect 138 13320 172 13354
rect 1666 13416 1700 13450
rect 138 13128 172 13162
rect 1666 13224 1700 13258
rect 138 12936 172 12970
rect 1666 13032 1700 13066
rect 138 12744 172 12778
rect 1666 12840 1700 12874
rect 138 12552 172 12586
rect 1666 12648 1700 12682
rect 138 12360 172 12394
rect 1666 12456 1700 12490
rect 138 12168 172 12202
rect 1666 12264 1700 12298
rect 138 11976 172 12010
rect 1666 12072 1700 12106
rect 138 11784 172 11818
rect 1666 11880 1700 11914
rect 138 11592 172 11626
rect 1666 11688 1700 11722
rect 138 11400 172 11434
rect 1666 11496 1700 11530
rect 138 11208 172 11242
rect 1666 11304 1700 11338
rect 138 11016 172 11050
rect 1666 11112 1700 11146
rect 138 10824 172 10858
rect 1666 10920 1700 10954
rect 138 10632 172 10666
rect 1666 10728 1700 10762
rect 138 10440 172 10474
rect 1666 10536 1700 10570
rect 138 10248 172 10282
rect 1666 10344 1700 10378
rect 138 10056 172 10090
rect 1666 10152 1700 10186
rect 138 9864 172 9898
rect 1666 9960 1700 9994
rect 138 9672 172 9706
rect 1666 9768 1700 9802
rect 138 9480 172 9514
rect 1666 9576 1700 9610
rect 138 9288 172 9322
rect 1666 9384 1700 9418
rect 138 9096 172 9130
rect 1666 9192 1700 9226
rect 138 8904 172 8938
rect 1666 9000 1700 9034
rect 138 8712 172 8746
rect 1666 8808 1700 8842
rect 138 8520 172 8554
rect 1666 8616 1700 8650
rect 138 8328 172 8362
rect 1666 8424 1700 8458
rect 138 8136 172 8170
rect 1666 8232 1700 8266
rect 138 7944 172 7978
rect 1666 8040 1700 8074
rect 138 7752 172 7786
rect 1666 7848 1700 7882
rect 138 7560 172 7594
rect 1666 7656 1700 7690
rect 138 7368 172 7402
rect 1666 7464 1700 7498
rect 138 7176 172 7210
rect 1666 7272 1700 7306
rect 138 6984 172 7018
rect 1666 7080 1700 7114
rect 138 6792 172 6826
rect 1666 6888 1700 6922
rect 138 6600 172 6634
rect 1666 6696 1700 6730
rect 138 6408 172 6442
rect 1666 6504 1700 6538
rect 138 6216 172 6250
rect 1666 6312 1700 6346
rect 138 6024 172 6058
rect 1666 6120 1700 6154
rect 138 5832 172 5866
rect 1666 5928 1700 5962
rect 138 5640 172 5674
rect 1666 5736 1700 5770
rect 138 5448 172 5482
rect 1666 5544 1700 5578
rect 138 5256 172 5290
rect 1666 5352 1700 5386
rect 138 5064 172 5098
rect 1666 5160 1700 5194
rect 138 4872 172 4906
rect 1666 4968 1700 5002
rect 138 4680 172 4714
rect 1666 4776 1700 4810
rect 138 4488 172 4522
rect 1666 4584 1700 4618
rect 138 4296 172 4330
rect 1666 4392 1700 4426
rect 138 4104 172 4138
rect 1666 4200 1700 4234
rect 138 3912 172 3946
rect 1666 4008 1700 4042
rect 138 3720 172 3754
rect 1666 3816 1700 3850
rect 138 3528 172 3562
rect 1666 3624 1700 3658
rect 138 3336 172 3370
rect 1666 3432 1700 3466
rect 138 3144 172 3178
rect 1666 3240 1700 3274
rect 138 2952 172 2986
rect 1666 3048 1700 3082
rect 138 2760 172 2794
rect 1666 2856 1700 2890
rect 138 2568 172 2602
rect 1666 2664 1700 2698
rect 138 2376 172 2410
rect 1666 2472 1700 2506
rect 138 2184 172 2218
rect 1666 2280 1700 2314
rect 138 1992 172 2026
rect 1666 2088 1700 2122
rect 138 1800 172 1834
rect 1666 1896 1700 1930
rect 138 1608 172 1642
rect 1666 1704 1700 1738
rect 138 1416 172 1450
rect 1666 1512 1700 1546
rect 138 1224 172 1258
rect 1666 1320 1700 1354
rect 138 1032 172 1066
rect 1666 1128 1700 1162
rect 138 840 172 874
rect 1666 936 1700 970
rect 1666 744 1700 778
<< locali >>
rect 36 21930 132 21964
rect 1706 21930 1802 21964
rect 36 21868 70 21930
rect 1768 21868 1802 21930
rect 138 21802 172 21818
rect 215 21816 231 21850
rect 1607 21816 1623 21850
rect 138 21752 172 21768
rect 215 21720 231 21754
rect 1607 21720 1623 21754
rect 1666 21706 1700 21722
rect 138 21610 172 21626
rect 215 21624 231 21658
rect 1607 21624 1623 21658
rect 1666 21656 1700 21672
rect 138 21560 172 21576
rect 215 21528 231 21562
rect 1607 21528 1623 21562
rect 1666 21514 1700 21530
rect 138 21418 172 21434
rect 215 21432 231 21466
rect 1607 21432 1623 21466
rect 1666 21464 1700 21480
rect 138 21368 172 21384
rect 215 21336 231 21370
rect 1607 21336 1623 21370
rect 1666 21322 1700 21338
rect 138 21226 172 21242
rect 215 21240 231 21274
rect 1607 21240 1623 21274
rect 1666 21272 1700 21288
rect 138 21176 172 21192
rect 215 21144 231 21178
rect 1607 21144 1623 21178
rect 1666 21130 1700 21146
rect 138 21034 172 21050
rect 215 21048 231 21082
rect 1607 21048 1623 21082
rect 1666 21080 1700 21096
rect 138 20984 172 21000
rect 215 20952 231 20986
rect 1607 20952 1623 20986
rect 1666 20938 1700 20954
rect 138 20842 172 20858
rect 215 20856 231 20890
rect 1607 20856 1623 20890
rect 1666 20888 1700 20904
rect 138 20792 172 20808
rect 215 20760 231 20794
rect 1607 20760 1623 20794
rect 1666 20746 1700 20762
rect 138 20650 172 20666
rect 215 20664 231 20698
rect 1607 20664 1623 20698
rect 1666 20696 1700 20712
rect 138 20600 172 20616
rect 215 20568 231 20602
rect 1607 20568 1623 20602
rect 1666 20554 1700 20570
rect 138 20458 172 20474
rect 215 20472 231 20506
rect 1607 20472 1623 20506
rect 1666 20504 1700 20520
rect 138 20408 172 20424
rect 215 20376 231 20410
rect 1607 20376 1623 20410
rect 1666 20362 1700 20378
rect 138 20266 172 20282
rect 215 20280 231 20314
rect 1607 20280 1623 20314
rect 1666 20312 1700 20328
rect 138 20216 172 20232
rect 215 20184 231 20218
rect 1607 20184 1623 20218
rect 1666 20170 1700 20186
rect 138 20074 172 20090
rect 215 20088 231 20122
rect 1607 20088 1623 20122
rect 1666 20120 1700 20136
rect 138 20024 172 20040
rect 215 19992 231 20026
rect 1607 19992 1623 20026
rect 1666 19978 1700 19994
rect 138 19882 172 19898
rect 215 19896 231 19930
rect 1607 19896 1623 19930
rect 1666 19928 1700 19944
rect 138 19832 172 19848
rect 215 19800 231 19834
rect 1607 19800 1623 19834
rect 1666 19786 1700 19802
rect 138 19690 172 19706
rect 215 19704 231 19738
rect 1607 19704 1623 19738
rect 1666 19736 1700 19752
rect 138 19640 172 19656
rect 215 19608 231 19642
rect 1607 19608 1623 19642
rect 1666 19594 1700 19610
rect 138 19498 172 19514
rect 215 19512 231 19546
rect 1607 19512 1623 19546
rect 1666 19544 1700 19560
rect 138 19448 172 19464
rect 215 19416 231 19450
rect 1607 19416 1623 19450
rect 1666 19402 1700 19418
rect 138 19306 172 19322
rect 215 19320 231 19354
rect 1607 19320 1623 19354
rect 1666 19352 1700 19368
rect 138 19256 172 19272
rect 215 19224 231 19258
rect 1607 19224 1623 19258
rect 1666 19210 1700 19226
rect 138 19114 172 19130
rect 215 19128 231 19162
rect 1607 19128 1623 19162
rect 1666 19160 1700 19176
rect 138 19064 172 19080
rect 215 19032 231 19066
rect 1607 19032 1623 19066
rect 1666 19018 1700 19034
rect 138 18922 172 18938
rect 215 18936 231 18970
rect 1607 18936 1623 18970
rect 1666 18968 1700 18984
rect 138 18872 172 18888
rect 215 18840 231 18874
rect 1607 18840 1623 18874
rect 1666 18826 1700 18842
rect 138 18730 172 18746
rect 215 18744 231 18778
rect 1607 18744 1623 18778
rect 1666 18776 1700 18792
rect 138 18680 172 18696
rect 215 18648 231 18682
rect 1607 18648 1623 18682
rect 1666 18634 1700 18650
rect 138 18538 172 18554
rect 215 18552 231 18586
rect 1607 18552 1623 18586
rect 1666 18584 1700 18600
rect 138 18488 172 18504
rect 215 18456 231 18490
rect 1607 18456 1623 18490
rect 1666 18442 1700 18458
rect 138 18346 172 18362
rect 215 18360 231 18394
rect 1607 18360 1623 18394
rect 1666 18392 1700 18408
rect 138 18296 172 18312
rect 215 18264 231 18298
rect 1607 18264 1623 18298
rect 1666 18250 1700 18266
rect 138 18154 172 18170
rect 215 18168 231 18202
rect 1607 18168 1623 18202
rect 1666 18200 1700 18216
rect 138 18104 172 18120
rect 215 18072 231 18106
rect 1607 18072 1623 18106
rect 1666 18058 1700 18074
rect 138 17962 172 17978
rect 215 17976 231 18010
rect 1607 17976 1623 18010
rect 1666 18008 1700 18024
rect 138 17912 172 17928
rect 215 17880 231 17914
rect 1607 17880 1623 17914
rect 1666 17866 1700 17882
rect 138 17770 172 17786
rect 215 17784 231 17818
rect 1607 17784 1623 17818
rect 1666 17816 1700 17832
rect 138 17720 172 17736
rect 215 17688 231 17722
rect 1607 17688 1623 17722
rect 1666 17674 1700 17690
rect 138 17578 172 17594
rect 215 17592 231 17626
rect 1607 17592 1623 17626
rect 1666 17624 1700 17640
rect 138 17528 172 17544
rect 215 17496 231 17530
rect 1607 17496 1623 17530
rect 1666 17482 1700 17498
rect 138 17386 172 17402
rect 215 17400 231 17434
rect 1607 17400 1623 17434
rect 1666 17432 1700 17448
rect 138 17336 172 17352
rect 215 17304 231 17338
rect 1607 17304 1623 17338
rect 1666 17290 1700 17306
rect 138 17194 172 17210
rect 215 17208 231 17242
rect 1607 17208 1623 17242
rect 1666 17240 1700 17256
rect 138 17144 172 17160
rect 215 17112 231 17146
rect 1607 17112 1623 17146
rect 1666 17098 1700 17114
rect 138 17002 172 17018
rect 215 17016 231 17050
rect 1607 17016 1623 17050
rect 1666 17048 1700 17064
rect 138 16952 172 16968
rect 215 16920 231 16954
rect 1607 16920 1623 16954
rect 1666 16906 1700 16922
rect 138 16810 172 16826
rect 215 16824 231 16858
rect 1607 16824 1623 16858
rect 1666 16856 1700 16872
rect 138 16760 172 16776
rect 215 16728 231 16762
rect 1607 16728 1623 16762
rect 1666 16714 1700 16730
rect 138 16618 172 16634
rect 215 16632 231 16666
rect 1607 16632 1623 16666
rect 1666 16664 1700 16680
rect 138 16568 172 16584
rect 215 16536 231 16570
rect 1607 16536 1623 16570
rect 1666 16522 1700 16538
rect 138 16426 172 16442
rect 215 16440 231 16474
rect 1607 16440 1623 16474
rect 1666 16472 1700 16488
rect 138 16376 172 16392
rect 215 16344 231 16378
rect 1607 16344 1623 16378
rect 1666 16330 1700 16346
rect 138 16234 172 16250
rect 215 16248 231 16282
rect 1607 16248 1623 16282
rect 1666 16280 1700 16296
rect 138 16184 172 16200
rect 215 16152 231 16186
rect 1607 16152 1623 16186
rect 1666 16138 1700 16154
rect 138 16042 172 16058
rect 215 16056 231 16090
rect 1607 16056 1623 16090
rect 1666 16088 1700 16104
rect 138 15992 172 16008
rect 215 15960 231 15994
rect 1607 15960 1623 15994
rect 1666 15946 1700 15962
rect 138 15850 172 15866
rect 215 15864 231 15898
rect 1607 15864 1623 15898
rect 1666 15896 1700 15912
rect 138 15800 172 15816
rect 215 15768 231 15802
rect 1607 15768 1623 15802
rect 1666 15754 1700 15770
rect 138 15658 172 15674
rect 215 15672 231 15706
rect 1607 15672 1623 15706
rect 1666 15704 1700 15720
rect 138 15608 172 15624
rect 215 15576 231 15610
rect 1607 15576 1623 15610
rect 1666 15562 1700 15578
rect 138 15466 172 15482
rect 215 15480 231 15514
rect 1607 15480 1623 15514
rect 1666 15512 1700 15528
rect 138 15416 172 15432
rect 215 15384 231 15418
rect 1607 15384 1623 15418
rect 1666 15370 1700 15386
rect 138 15274 172 15290
rect 215 15288 231 15322
rect 1607 15288 1623 15322
rect 1666 15320 1700 15336
rect 138 15224 172 15240
rect 215 15192 231 15226
rect 1607 15192 1623 15226
rect 1666 15178 1700 15194
rect 138 15082 172 15098
rect 215 15096 231 15130
rect 1607 15096 1623 15130
rect 1666 15128 1700 15144
rect 138 15032 172 15048
rect 215 15000 231 15034
rect 1607 15000 1623 15034
rect 1666 14986 1700 15002
rect 138 14890 172 14906
rect 215 14904 231 14938
rect 1607 14904 1623 14938
rect 1666 14936 1700 14952
rect 138 14840 172 14856
rect 215 14808 231 14842
rect 1607 14808 1623 14842
rect 1666 14794 1700 14810
rect 138 14698 172 14714
rect 215 14712 231 14746
rect 1607 14712 1623 14746
rect 1666 14744 1700 14760
rect 138 14648 172 14664
rect 215 14616 231 14650
rect 1607 14616 1623 14650
rect 1666 14602 1700 14618
rect 138 14506 172 14522
rect 215 14520 231 14554
rect 1607 14520 1623 14554
rect 1666 14552 1700 14568
rect 138 14456 172 14472
rect 215 14424 231 14458
rect 1607 14424 1623 14458
rect 1666 14410 1700 14426
rect 138 14314 172 14330
rect 215 14328 231 14362
rect 1607 14328 1623 14362
rect 1666 14360 1700 14376
rect 138 14264 172 14280
rect 215 14232 231 14266
rect 1607 14232 1623 14266
rect 1666 14218 1700 14234
rect 138 14122 172 14138
rect 215 14136 231 14170
rect 1607 14136 1623 14170
rect 1666 14168 1700 14184
rect 138 14072 172 14088
rect 215 14040 231 14074
rect 1607 14040 1623 14074
rect 1666 14026 1700 14042
rect 138 13930 172 13946
rect 215 13944 231 13978
rect 1607 13944 1623 13978
rect 1666 13976 1700 13992
rect 138 13880 172 13896
rect 215 13848 231 13882
rect 1607 13848 1623 13882
rect 1666 13834 1700 13850
rect 138 13738 172 13754
rect 215 13752 231 13786
rect 1607 13752 1623 13786
rect 1666 13784 1700 13800
rect 138 13688 172 13704
rect 215 13656 231 13690
rect 1607 13656 1623 13690
rect 1666 13642 1700 13658
rect 138 13546 172 13562
rect 215 13560 231 13594
rect 1607 13560 1623 13594
rect 1666 13592 1700 13608
rect 138 13496 172 13512
rect 215 13464 231 13498
rect 1607 13464 1623 13498
rect 1666 13450 1700 13466
rect 138 13354 172 13370
rect 215 13368 231 13402
rect 1607 13368 1623 13402
rect 1666 13400 1700 13416
rect 138 13304 172 13320
rect 215 13272 231 13306
rect 1607 13272 1623 13306
rect 1666 13258 1700 13274
rect 138 13162 172 13178
rect 215 13176 231 13210
rect 1607 13176 1623 13210
rect 1666 13208 1700 13224
rect 138 13112 172 13128
rect 215 13080 231 13114
rect 1607 13080 1623 13114
rect 1666 13066 1700 13082
rect 138 12970 172 12986
rect 215 12984 231 13018
rect 1607 12984 1623 13018
rect 1666 13016 1700 13032
rect 138 12920 172 12936
rect 215 12888 231 12922
rect 1607 12888 1623 12922
rect 1666 12874 1700 12890
rect 138 12778 172 12794
rect 215 12792 231 12826
rect 1607 12792 1623 12826
rect 1666 12824 1700 12840
rect 138 12728 172 12744
rect 215 12696 231 12730
rect 1607 12696 1623 12730
rect 1666 12682 1700 12698
rect 138 12586 172 12602
rect 215 12600 231 12634
rect 1607 12600 1623 12634
rect 1666 12632 1700 12648
rect 138 12536 172 12552
rect 215 12504 231 12538
rect 1607 12504 1623 12538
rect 1666 12490 1700 12506
rect 138 12394 172 12410
rect 215 12408 231 12442
rect 1607 12408 1623 12442
rect 1666 12440 1700 12456
rect 138 12344 172 12360
rect 215 12312 231 12346
rect 1607 12312 1623 12346
rect 1666 12298 1700 12314
rect 138 12202 172 12218
rect 215 12216 231 12250
rect 1607 12216 1623 12250
rect 1666 12248 1700 12264
rect 138 12152 172 12168
rect 215 12120 231 12154
rect 1607 12120 1623 12154
rect 1666 12106 1700 12122
rect 138 12010 172 12026
rect 215 12024 231 12058
rect 1607 12024 1623 12058
rect 1666 12056 1700 12072
rect 138 11960 172 11976
rect 215 11928 231 11962
rect 1607 11928 1623 11962
rect 1666 11914 1700 11930
rect 138 11818 172 11834
rect 215 11832 231 11866
rect 1607 11832 1623 11866
rect 1666 11864 1700 11880
rect 138 11768 172 11784
rect 215 11736 231 11770
rect 1607 11736 1623 11770
rect 1666 11722 1700 11738
rect 138 11626 172 11642
rect 215 11640 231 11674
rect 1607 11640 1623 11674
rect 1666 11672 1700 11688
rect 138 11576 172 11592
rect 215 11544 231 11578
rect 1607 11544 1623 11578
rect 1666 11530 1700 11546
rect 138 11434 172 11450
rect 215 11448 231 11482
rect 1607 11448 1623 11482
rect 1666 11480 1700 11496
rect 138 11384 172 11400
rect 215 11352 231 11386
rect 1607 11352 1623 11386
rect 1666 11338 1700 11354
rect 138 11242 172 11258
rect 215 11256 231 11290
rect 1607 11256 1623 11290
rect 1666 11288 1700 11304
rect 138 11192 172 11208
rect 215 11160 231 11194
rect 1607 11160 1623 11194
rect 1666 11146 1700 11162
rect 138 11050 172 11066
rect 215 11064 231 11098
rect 1607 11064 1623 11098
rect 1666 11096 1700 11112
rect 138 11000 172 11016
rect 215 10968 231 11002
rect 1607 10968 1623 11002
rect 1666 10954 1700 10970
rect 138 10858 172 10874
rect 215 10872 231 10906
rect 1607 10872 1623 10906
rect 1666 10904 1700 10920
rect 138 10808 172 10824
rect 215 10776 231 10810
rect 1607 10776 1623 10810
rect 1666 10762 1700 10778
rect 138 10666 172 10682
rect 215 10680 231 10714
rect 1607 10680 1623 10714
rect 1666 10712 1700 10728
rect 138 10616 172 10632
rect 215 10584 231 10618
rect 1607 10584 1623 10618
rect 1666 10570 1700 10586
rect 138 10474 172 10490
rect 215 10488 231 10522
rect 1607 10488 1623 10522
rect 1666 10520 1700 10536
rect 138 10424 172 10440
rect 215 10392 231 10426
rect 1607 10392 1623 10426
rect 1666 10378 1700 10394
rect 138 10282 172 10298
rect 215 10296 231 10330
rect 1607 10296 1623 10330
rect 1666 10328 1700 10344
rect 138 10232 172 10248
rect 215 10200 231 10234
rect 1607 10200 1623 10234
rect 1666 10186 1700 10202
rect 138 10090 172 10106
rect 215 10104 231 10138
rect 1607 10104 1623 10138
rect 1666 10136 1700 10152
rect 138 10040 172 10056
rect 215 10008 231 10042
rect 1607 10008 1623 10042
rect 1666 9994 1700 10010
rect 138 9898 172 9914
rect 215 9912 231 9946
rect 1607 9912 1623 9946
rect 1666 9944 1700 9960
rect 138 9848 172 9864
rect 215 9816 231 9850
rect 1607 9816 1623 9850
rect 1666 9802 1700 9818
rect 138 9706 172 9722
rect 215 9720 231 9754
rect 1607 9720 1623 9754
rect 1666 9752 1700 9768
rect 138 9656 172 9672
rect 215 9624 231 9658
rect 1607 9624 1623 9658
rect 1666 9610 1700 9626
rect 138 9514 172 9530
rect 215 9528 231 9562
rect 1607 9528 1623 9562
rect 1666 9560 1700 9576
rect 138 9464 172 9480
rect 215 9432 231 9466
rect 1607 9432 1623 9466
rect 1666 9418 1700 9434
rect 138 9322 172 9338
rect 215 9336 231 9370
rect 1607 9336 1623 9370
rect 1666 9368 1700 9384
rect 138 9272 172 9288
rect 215 9240 231 9274
rect 1607 9240 1623 9274
rect 1666 9226 1700 9242
rect 138 9130 172 9146
rect 215 9144 231 9178
rect 1607 9144 1623 9178
rect 1666 9176 1700 9192
rect 138 9080 172 9096
rect 215 9048 231 9082
rect 1607 9048 1623 9082
rect 1666 9034 1700 9050
rect 138 8938 172 8954
rect 215 8952 231 8986
rect 1607 8952 1623 8986
rect 1666 8984 1700 9000
rect 138 8888 172 8904
rect 215 8856 231 8890
rect 1607 8856 1623 8890
rect 1666 8842 1700 8858
rect 138 8746 172 8762
rect 215 8760 231 8794
rect 1607 8760 1623 8794
rect 1666 8792 1700 8808
rect 138 8696 172 8712
rect 215 8664 231 8698
rect 1607 8664 1623 8698
rect 1666 8650 1700 8666
rect 138 8554 172 8570
rect 215 8568 231 8602
rect 1607 8568 1623 8602
rect 1666 8600 1700 8616
rect 138 8504 172 8520
rect 215 8472 231 8506
rect 1607 8472 1623 8506
rect 1666 8458 1700 8474
rect 138 8362 172 8378
rect 215 8376 231 8410
rect 1607 8376 1623 8410
rect 1666 8408 1700 8424
rect 138 8312 172 8328
rect 215 8280 231 8314
rect 1607 8280 1623 8314
rect 1666 8266 1700 8282
rect 138 8170 172 8186
rect 215 8184 231 8218
rect 1607 8184 1623 8218
rect 1666 8216 1700 8232
rect 138 8120 172 8136
rect 215 8088 231 8122
rect 1607 8088 1623 8122
rect 1666 8074 1700 8090
rect 138 7978 172 7994
rect 215 7992 231 8026
rect 1607 7992 1623 8026
rect 1666 8024 1700 8040
rect 138 7928 172 7944
rect 215 7896 231 7930
rect 1607 7896 1623 7930
rect 1666 7882 1700 7898
rect 138 7786 172 7802
rect 215 7800 231 7834
rect 1607 7800 1623 7834
rect 1666 7832 1700 7848
rect 138 7736 172 7752
rect 215 7704 231 7738
rect 1607 7704 1623 7738
rect 1666 7690 1700 7706
rect 138 7594 172 7610
rect 215 7608 231 7642
rect 1607 7608 1623 7642
rect 1666 7640 1700 7656
rect 138 7544 172 7560
rect 215 7512 231 7546
rect 1607 7512 1623 7546
rect 1666 7498 1700 7514
rect 138 7402 172 7418
rect 215 7416 231 7450
rect 1607 7416 1623 7450
rect 1666 7448 1700 7464
rect 138 7352 172 7368
rect 215 7320 231 7354
rect 1607 7320 1623 7354
rect 1666 7306 1700 7322
rect 138 7210 172 7226
rect 215 7224 231 7258
rect 1607 7224 1623 7258
rect 1666 7256 1700 7272
rect 138 7160 172 7176
rect 215 7128 231 7162
rect 1607 7128 1623 7162
rect 1666 7114 1700 7130
rect 138 7018 172 7034
rect 215 7032 231 7066
rect 1607 7032 1623 7066
rect 1666 7064 1700 7080
rect 138 6968 172 6984
rect 215 6936 231 6970
rect 1607 6936 1623 6970
rect 1666 6922 1700 6938
rect 138 6826 172 6842
rect 215 6840 231 6874
rect 1607 6840 1623 6874
rect 1666 6872 1700 6888
rect 138 6776 172 6792
rect 215 6744 231 6778
rect 1607 6744 1623 6778
rect 1666 6730 1700 6746
rect 138 6634 172 6650
rect 215 6648 231 6682
rect 1607 6648 1623 6682
rect 1666 6680 1700 6696
rect 138 6584 172 6600
rect 215 6552 231 6586
rect 1607 6552 1623 6586
rect 1666 6538 1700 6554
rect 138 6442 172 6458
rect 215 6456 231 6490
rect 1607 6456 1623 6490
rect 1666 6488 1700 6504
rect 138 6392 172 6408
rect 215 6360 231 6394
rect 1607 6360 1623 6394
rect 1666 6346 1700 6362
rect 138 6250 172 6266
rect 215 6264 231 6298
rect 1607 6264 1623 6298
rect 1666 6296 1700 6312
rect 138 6200 172 6216
rect 215 6168 231 6202
rect 1607 6168 1623 6202
rect 1666 6154 1700 6170
rect 138 6058 172 6074
rect 215 6072 231 6106
rect 1607 6072 1623 6106
rect 1666 6104 1700 6120
rect 138 6008 172 6024
rect 215 5976 231 6010
rect 1607 5976 1623 6010
rect 1666 5962 1700 5978
rect 138 5866 172 5882
rect 215 5880 231 5914
rect 1607 5880 1623 5914
rect 1666 5912 1700 5928
rect 138 5816 172 5832
rect 215 5784 231 5818
rect 1607 5784 1623 5818
rect 1666 5770 1700 5786
rect 138 5674 172 5690
rect 215 5688 231 5722
rect 1607 5688 1623 5722
rect 1666 5720 1700 5736
rect 138 5624 172 5640
rect 215 5592 231 5626
rect 1607 5592 1623 5626
rect 1666 5578 1700 5594
rect 138 5482 172 5498
rect 215 5496 231 5530
rect 1607 5496 1623 5530
rect 1666 5528 1700 5544
rect 138 5432 172 5448
rect 215 5400 231 5434
rect 1607 5400 1623 5434
rect 1666 5386 1700 5402
rect 138 5290 172 5306
rect 215 5304 231 5338
rect 1607 5304 1623 5338
rect 1666 5336 1700 5352
rect 138 5240 172 5256
rect 215 5208 231 5242
rect 1607 5208 1623 5242
rect 1666 5194 1700 5210
rect 138 5098 172 5114
rect 215 5112 231 5146
rect 1607 5112 1623 5146
rect 1666 5144 1700 5160
rect 138 5048 172 5064
rect 215 5016 231 5050
rect 1607 5016 1623 5050
rect 1666 5002 1700 5018
rect 138 4906 172 4922
rect 215 4920 231 4954
rect 1607 4920 1623 4954
rect 1666 4952 1700 4968
rect 138 4856 172 4872
rect 215 4824 231 4858
rect 1607 4824 1623 4858
rect 1666 4810 1700 4826
rect 138 4714 172 4730
rect 215 4728 231 4762
rect 1607 4728 1623 4762
rect 1666 4760 1700 4776
rect 138 4664 172 4680
rect 215 4632 231 4666
rect 1607 4632 1623 4666
rect 1666 4618 1700 4634
rect 138 4522 172 4538
rect 215 4536 231 4570
rect 1607 4536 1623 4570
rect 1666 4568 1700 4584
rect 138 4472 172 4488
rect 215 4440 231 4474
rect 1607 4440 1623 4474
rect 1666 4426 1700 4442
rect 138 4330 172 4346
rect 215 4344 231 4378
rect 1607 4344 1623 4378
rect 1666 4376 1700 4392
rect 138 4280 172 4296
rect 215 4248 231 4282
rect 1607 4248 1623 4282
rect 1666 4234 1700 4250
rect 138 4138 172 4154
rect 215 4152 231 4186
rect 1607 4152 1623 4186
rect 1666 4184 1700 4200
rect 138 4088 172 4104
rect 215 4056 231 4090
rect 1607 4056 1623 4090
rect 1666 4042 1700 4058
rect 138 3946 172 3962
rect 215 3960 231 3994
rect 1607 3960 1623 3994
rect 1666 3992 1700 4008
rect 138 3896 172 3912
rect 215 3864 231 3898
rect 1607 3864 1623 3898
rect 1666 3850 1700 3866
rect 138 3754 172 3770
rect 215 3768 231 3802
rect 1607 3768 1623 3802
rect 1666 3800 1700 3816
rect 138 3704 172 3720
rect 215 3672 231 3706
rect 1607 3672 1623 3706
rect 1666 3658 1700 3674
rect 138 3562 172 3578
rect 215 3576 231 3610
rect 1607 3576 1623 3610
rect 1666 3608 1700 3624
rect 138 3512 172 3528
rect 215 3480 231 3514
rect 1607 3480 1623 3514
rect 1666 3466 1700 3482
rect 138 3370 172 3386
rect 215 3384 231 3418
rect 1607 3384 1623 3418
rect 1666 3416 1700 3432
rect 138 3320 172 3336
rect 215 3288 231 3322
rect 1607 3288 1623 3322
rect 1666 3274 1700 3290
rect 138 3178 172 3194
rect 215 3192 231 3226
rect 1607 3192 1623 3226
rect 1666 3224 1700 3240
rect 138 3128 172 3144
rect 215 3096 231 3130
rect 1607 3096 1623 3130
rect 1666 3082 1700 3098
rect 138 2986 172 3002
rect 215 3000 231 3034
rect 1607 3000 1623 3034
rect 1666 3032 1700 3048
rect 138 2936 172 2952
rect 215 2904 231 2938
rect 1607 2904 1623 2938
rect 1666 2890 1700 2906
rect 138 2794 172 2810
rect 215 2808 231 2842
rect 1607 2808 1623 2842
rect 1666 2840 1700 2856
rect 138 2744 172 2760
rect 215 2712 231 2746
rect 1607 2712 1623 2746
rect 1666 2698 1700 2714
rect 138 2602 172 2618
rect 215 2616 231 2650
rect 1607 2616 1623 2650
rect 1666 2648 1700 2664
rect 138 2552 172 2568
rect 215 2520 231 2554
rect 1607 2520 1623 2554
rect 1666 2506 1700 2522
rect 138 2410 172 2426
rect 215 2424 231 2458
rect 1607 2424 1623 2458
rect 1666 2456 1700 2472
rect 138 2360 172 2376
rect 215 2328 231 2362
rect 1607 2328 1623 2362
rect 1666 2314 1700 2330
rect 138 2218 172 2234
rect 215 2232 231 2266
rect 1607 2232 1623 2266
rect 1666 2264 1700 2280
rect 138 2168 172 2184
rect 215 2136 231 2170
rect 1607 2136 1623 2170
rect 1666 2122 1700 2138
rect 138 2026 172 2042
rect 215 2040 231 2074
rect 1607 2040 1623 2074
rect 1666 2072 1700 2088
rect 138 1976 172 1992
rect 215 1944 231 1978
rect 1607 1944 1623 1978
rect 1666 1930 1700 1946
rect 138 1834 172 1850
rect 215 1848 231 1882
rect 1607 1848 1623 1882
rect 1666 1880 1700 1896
rect 138 1784 172 1800
rect 215 1752 231 1786
rect 1607 1752 1623 1786
rect 1666 1738 1700 1754
rect 138 1642 172 1658
rect 215 1656 231 1690
rect 1607 1656 1623 1690
rect 1666 1688 1700 1704
rect 138 1592 172 1608
rect 215 1560 231 1594
rect 1607 1560 1623 1594
rect 1666 1546 1700 1562
rect 138 1450 172 1466
rect 215 1464 231 1498
rect 1607 1464 1623 1498
rect 1666 1496 1700 1512
rect 138 1400 172 1416
rect 215 1368 231 1402
rect 1607 1368 1623 1402
rect 1666 1354 1700 1370
rect 138 1258 172 1274
rect 215 1272 231 1306
rect 1607 1272 1623 1306
rect 1666 1304 1700 1320
rect 138 1208 172 1224
rect 215 1176 231 1210
rect 1607 1176 1623 1210
rect 1666 1162 1700 1178
rect 138 1066 172 1082
rect 215 1080 231 1114
rect 1607 1080 1623 1114
rect 1666 1112 1700 1128
rect 138 1016 172 1032
rect 215 984 231 1018
rect 1607 984 1623 1018
rect 1666 970 1700 986
rect 138 874 172 890
rect 215 888 231 922
rect 1607 888 1623 922
rect 1666 920 1700 936
rect 138 824 172 840
rect 215 792 231 826
rect 1607 792 1623 826
rect 1666 778 1700 794
rect 215 696 231 730
rect 1607 696 1623 730
rect 1666 728 1700 744
rect 36 616 70 678
rect 1768 616 1802 678
rect 36 582 132 616
rect 1706 582 1802 616
<< viali >>
rect 231 21816 1607 21850
rect 138 21768 172 21802
rect 231 21720 1607 21754
rect 1666 21672 1700 21706
rect 231 21624 1607 21658
rect 138 21576 172 21610
rect 231 21528 1607 21562
rect 1666 21480 1700 21514
rect 231 21432 1607 21466
rect 138 21384 172 21418
rect 231 21336 1607 21370
rect 1666 21288 1700 21322
rect 231 21240 1607 21274
rect 138 21192 172 21226
rect 231 21144 1607 21178
rect 1666 21096 1700 21130
rect 231 21048 1607 21082
rect 138 21000 172 21034
rect 231 20952 1607 20986
rect 1666 20904 1700 20938
rect 231 20856 1607 20890
rect 138 20808 172 20842
rect 231 20760 1607 20794
rect 1666 20712 1700 20746
rect 231 20664 1607 20698
rect 138 20616 172 20650
rect 231 20568 1607 20602
rect 1666 20520 1700 20554
rect 231 20472 1607 20506
rect 138 20424 172 20458
rect 231 20376 1607 20410
rect 1666 20328 1700 20362
rect 231 20280 1607 20314
rect 138 20232 172 20266
rect 231 20184 1607 20218
rect 1666 20136 1700 20170
rect 231 20088 1607 20122
rect 138 20040 172 20074
rect 231 19992 1607 20026
rect 1666 19944 1700 19978
rect 231 19896 1607 19930
rect 138 19848 172 19882
rect 231 19800 1607 19834
rect 1666 19752 1700 19786
rect 231 19704 1607 19738
rect 138 19656 172 19690
rect 231 19608 1607 19642
rect 1666 19560 1700 19594
rect 231 19512 1607 19546
rect 138 19464 172 19498
rect 231 19416 1607 19450
rect 1666 19368 1700 19402
rect 231 19320 1607 19354
rect 138 19272 172 19306
rect 231 19224 1607 19258
rect 1666 19176 1700 19210
rect 231 19128 1607 19162
rect 138 19080 172 19114
rect 231 19032 1607 19066
rect 1666 18984 1700 19018
rect 231 18936 1607 18970
rect 138 18888 172 18922
rect 231 18840 1607 18874
rect 1666 18792 1700 18826
rect 231 18744 1607 18778
rect 138 18696 172 18730
rect 231 18648 1607 18682
rect 1666 18600 1700 18634
rect 231 18552 1607 18586
rect 138 18504 172 18538
rect 231 18456 1607 18490
rect 1666 18408 1700 18442
rect 231 18360 1607 18394
rect 138 18312 172 18346
rect 231 18264 1607 18298
rect 1666 18216 1700 18250
rect 231 18168 1607 18202
rect 138 18120 172 18154
rect 231 18072 1607 18106
rect 1666 18024 1700 18058
rect 231 17976 1607 18010
rect 138 17928 172 17962
rect 231 17880 1607 17914
rect 1666 17832 1700 17866
rect 231 17784 1607 17818
rect 138 17736 172 17770
rect 231 17688 1607 17722
rect 1666 17640 1700 17674
rect 231 17592 1607 17626
rect 138 17544 172 17578
rect 231 17496 1607 17530
rect 1666 17448 1700 17482
rect 231 17400 1607 17434
rect 138 17352 172 17386
rect 231 17304 1607 17338
rect 1666 17256 1700 17290
rect 231 17208 1607 17242
rect 138 17160 172 17194
rect 231 17112 1607 17146
rect 1666 17064 1700 17098
rect 231 17016 1607 17050
rect 138 16968 172 17002
rect 231 16920 1607 16954
rect 1666 16872 1700 16906
rect 231 16824 1607 16858
rect 138 16776 172 16810
rect 231 16728 1607 16762
rect 1666 16680 1700 16714
rect 231 16632 1607 16666
rect 138 16584 172 16618
rect 231 16536 1607 16570
rect 1666 16488 1700 16522
rect 231 16440 1607 16474
rect 138 16392 172 16426
rect 231 16344 1607 16378
rect 1666 16296 1700 16330
rect 231 16248 1607 16282
rect 138 16200 172 16234
rect 231 16152 1607 16186
rect 1666 16104 1700 16138
rect 231 16056 1607 16090
rect 138 16008 172 16042
rect 231 15960 1607 15994
rect 1666 15912 1700 15946
rect 231 15864 1607 15898
rect 138 15816 172 15850
rect 231 15768 1607 15802
rect 1666 15720 1700 15754
rect 231 15672 1607 15706
rect 138 15624 172 15658
rect 231 15576 1607 15610
rect 1666 15528 1700 15562
rect 231 15480 1607 15514
rect 138 15432 172 15466
rect 231 15384 1607 15418
rect 1666 15336 1700 15370
rect 231 15288 1607 15322
rect 138 15240 172 15274
rect 231 15192 1607 15226
rect 1666 15144 1700 15178
rect 231 15096 1607 15130
rect 138 15048 172 15082
rect 231 15000 1607 15034
rect 1666 14952 1700 14986
rect 231 14904 1607 14938
rect 138 14856 172 14890
rect 231 14808 1607 14842
rect 1666 14760 1700 14794
rect 231 14712 1607 14746
rect 138 14664 172 14698
rect 231 14616 1607 14650
rect 1666 14568 1700 14602
rect 231 14520 1607 14554
rect 138 14472 172 14506
rect 231 14424 1607 14458
rect 1666 14376 1700 14410
rect 231 14328 1607 14362
rect 138 14280 172 14314
rect 231 14232 1607 14266
rect 1666 14184 1700 14218
rect 231 14136 1607 14170
rect 138 14088 172 14122
rect 231 14040 1607 14074
rect 1666 13992 1700 14026
rect 231 13944 1607 13978
rect 138 13896 172 13930
rect 231 13848 1607 13882
rect 1666 13800 1700 13834
rect 231 13752 1607 13786
rect 138 13704 172 13738
rect 231 13656 1607 13690
rect 1666 13608 1700 13642
rect 231 13560 1607 13594
rect 138 13512 172 13546
rect 231 13464 1607 13498
rect 1666 13416 1700 13450
rect 231 13368 1607 13402
rect 138 13320 172 13354
rect 231 13272 1607 13306
rect 1666 13224 1700 13258
rect 231 13176 1607 13210
rect 138 13128 172 13162
rect 231 13080 1607 13114
rect 1666 13032 1700 13066
rect 231 12984 1607 13018
rect 138 12936 172 12970
rect 231 12888 1607 12922
rect 1666 12840 1700 12874
rect 231 12792 1607 12826
rect 138 12744 172 12778
rect 231 12696 1607 12730
rect 1666 12648 1700 12682
rect 231 12600 1607 12634
rect 138 12552 172 12586
rect 231 12504 1607 12538
rect 1666 12456 1700 12490
rect 231 12408 1607 12442
rect 138 12360 172 12394
rect 231 12312 1607 12346
rect 1666 12264 1700 12298
rect 231 12216 1607 12250
rect 138 12168 172 12202
rect 231 12120 1607 12154
rect 1666 12072 1700 12106
rect 231 12024 1607 12058
rect 138 11976 172 12010
rect 231 11928 1607 11962
rect 1666 11880 1700 11914
rect 231 11832 1607 11866
rect 138 11784 172 11818
rect 231 11736 1607 11770
rect 1666 11688 1700 11722
rect 231 11640 1607 11674
rect 138 11592 172 11626
rect 231 11544 1607 11578
rect 1666 11496 1700 11530
rect 231 11448 1607 11482
rect 138 11400 172 11434
rect 231 11352 1607 11386
rect 1666 11304 1700 11338
rect 231 11256 1607 11290
rect 138 11208 172 11242
rect 231 11160 1607 11194
rect 1666 11112 1700 11146
rect 231 11064 1607 11098
rect 138 11016 172 11050
rect 231 10968 1607 11002
rect 1666 10920 1700 10954
rect 231 10872 1607 10906
rect 138 10824 172 10858
rect 231 10776 1607 10810
rect 1666 10728 1700 10762
rect 231 10680 1607 10714
rect 138 10632 172 10666
rect 231 10584 1607 10618
rect 1666 10536 1700 10570
rect 231 10488 1607 10522
rect 138 10440 172 10474
rect 231 10392 1607 10426
rect 1666 10344 1700 10378
rect 231 10296 1607 10330
rect 138 10248 172 10282
rect 231 10200 1607 10234
rect 1666 10152 1700 10186
rect 231 10104 1607 10138
rect 138 10056 172 10090
rect 231 10008 1607 10042
rect 1666 9960 1700 9994
rect 231 9912 1607 9946
rect 138 9864 172 9898
rect 231 9816 1607 9850
rect 1666 9768 1700 9802
rect 231 9720 1607 9754
rect 138 9672 172 9706
rect 231 9624 1607 9658
rect 1666 9576 1700 9610
rect 231 9528 1607 9562
rect 138 9480 172 9514
rect 231 9432 1607 9466
rect 1666 9384 1700 9418
rect 231 9336 1607 9370
rect 138 9288 172 9322
rect 231 9240 1607 9274
rect 1666 9192 1700 9226
rect 231 9144 1607 9178
rect 138 9096 172 9130
rect 231 9048 1607 9082
rect 1666 9000 1700 9034
rect 231 8952 1607 8986
rect 138 8904 172 8938
rect 231 8856 1607 8890
rect 1666 8808 1700 8842
rect 231 8760 1607 8794
rect 138 8712 172 8746
rect 231 8664 1607 8698
rect 1666 8616 1700 8650
rect 231 8568 1607 8602
rect 138 8520 172 8554
rect 231 8472 1607 8506
rect 1666 8424 1700 8458
rect 231 8376 1607 8410
rect 138 8328 172 8362
rect 231 8280 1607 8314
rect 1666 8232 1700 8266
rect 231 8184 1607 8218
rect 138 8136 172 8170
rect 231 8088 1607 8122
rect 1666 8040 1700 8074
rect 231 7992 1607 8026
rect 138 7944 172 7978
rect 231 7896 1607 7930
rect 1666 7848 1700 7882
rect 231 7800 1607 7834
rect 138 7752 172 7786
rect 231 7704 1607 7738
rect 1666 7656 1700 7690
rect 231 7608 1607 7642
rect 138 7560 172 7594
rect 231 7512 1607 7546
rect 1666 7464 1700 7498
rect 231 7416 1607 7450
rect 138 7368 172 7402
rect 231 7320 1607 7354
rect 1666 7272 1700 7306
rect 231 7224 1607 7258
rect 138 7176 172 7210
rect 231 7128 1607 7162
rect 1666 7080 1700 7114
rect 231 7032 1607 7066
rect 138 6984 172 7018
rect 231 6936 1607 6970
rect 1666 6888 1700 6922
rect 231 6840 1607 6874
rect 138 6792 172 6826
rect 231 6744 1607 6778
rect 1666 6696 1700 6730
rect 231 6648 1607 6682
rect 138 6600 172 6634
rect 231 6552 1607 6586
rect 1666 6504 1700 6538
rect 231 6456 1607 6490
rect 138 6408 172 6442
rect 231 6360 1607 6394
rect 1666 6312 1700 6346
rect 231 6264 1607 6298
rect 138 6216 172 6250
rect 231 6168 1607 6202
rect 1666 6120 1700 6154
rect 231 6072 1607 6106
rect 138 6024 172 6058
rect 231 5976 1607 6010
rect 1666 5928 1700 5962
rect 231 5880 1607 5914
rect 138 5832 172 5866
rect 231 5784 1607 5818
rect 1666 5736 1700 5770
rect 231 5688 1607 5722
rect 138 5640 172 5674
rect 231 5592 1607 5626
rect 1666 5544 1700 5578
rect 231 5496 1607 5530
rect 138 5448 172 5482
rect 231 5400 1607 5434
rect 1666 5352 1700 5386
rect 231 5304 1607 5338
rect 138 5256 172 5290
rect 231 5208 1607 5242
rect 1666 5160 1700 5194
rect 231 5112 1607 5146
rect 138 5064 172 5098
rect 231 5016 1607 5050
rect 1666 4968 1700 5002
rect 231 4920 1607 4954
rect 138 4872 172 4906
rect 231 4824 1607 4858
rect 1666 4776 1700 4810
rect 231 4728 1607 4762
rect 138 4680 172 4714
rect 231 4632 1607 4666
rect 1666 4584 1700 4618
rect 231 4536 1607 4570
rect 138 4488 172 4522
rect 231 4440 1607 4474
rect 1666 4392 1700 4426
rect 231 4344 1607 4378
rect 138 4296 172 4330
rect 231 4248 1607 4282
rect 1666 4200 1700 4234
rect 231 4152 1607 4186
rect 138 4104 172 4138
rect 231 4056 1607 4090
rect 1666 4008 1700 4042
rect 231 3960 1607 3994
rect 138 3912 172 3946
rect 231 3864 1607 3898
rect 1666 3816 1700 3850
rect 231 3768 1607 3802
rect 138 3720 172 3754
rect 231 3672 1607 3706
rect 1666 3624 1700 3658
rect 231 3576 1607 3610
rect 138 3528 172 3562
rect 231 3480 1607 3514
rect 1666 3432 1700 3466
rect 231 3384 1607 3418
rect 138 3336 172 3370
rect 231 3288 1607 3322
rect 1666 3240 1700 3274
rect 231 3192 1607 3226
rect 138 3144 172 3178
rect 231 3096 1607 3130
rect 1666 3048 1700 3082
rect 231 3000 1607 3034
rect 138 2952 172 2986
rect 231 2904 1607 2938
rect 1666 2856 1700 2890
rect 231 2808 1607 2842
rect 138 2760 172 2794
rect 231 2712 1607 2746
rect 1666 2664 1700 2698
rect 231 2616 1607 2650
rect 138 2568 172 2602
rect 231 2520 1607 2554
rect 1666 2472 1700 2506
rect 231 2424 1607 2458
rect 138 2376 172 2410
rect 231 2328 1607 2362
rect 1666 2280 1700 2314
rect 231 2232 1607 2266
rect 138 2184 172 2218
rect 231 2136 1607 2170
rect 1666 2088 1700 2122
rect 231 2040 1607 2074
rect 138 1992 172 2026
rect 231 1944 1607 1978
rect 1666 1896 1700 1930
rect 231 1848 1607 1882
rect 138 1800 172 1834
rect 231 1752 1607 1786
rect 1666 1704 1700 1738
rect 231 1656 1607 1690
rect 138 1608 172 1642
rect 231 1560 1607 1594
rect 1666 1512 1700 1546
rect 231 1464 1607 1498
rect 138 1416 172 1450
rect 231 1368 1607 1402
rect 1666 1320 1700 1354
rect 231 1272 1607 1306
rect 138 1224 172 1258
rect 231 1176 1607 1210
rect 1666 1128 1700 1162
rect 231 1080 1607 1114
rect 138 1032 172 1066
rect 231 984 1607 1018
rect 1666 936 1700 970
rect 231 888 1607 922
rect 138 840 172 874
rect 231 792 1607 826
rect 1666 744 1700 778
rect 231 696 1607 730
<< metal1 >>
rect 219 21850 1619 21856
rect 219 21816 231 21850
rect 1607 21816 1619 21850
rect 132 21802 178 21814
rect 219 21810 1619 21816
rect 132 21768 138 21802
rect 172 21768 178 21802
rect 132 21756 178 21768
rect 219 21754 1619 21760
rect 219 21720 231 21754
rect 1607 21720 1619 21754
rect 219 21714 1619 21720
rect 1660 21706 1706 21718
rect 1660 21672 1666 21706
rect 1700 21672 1706 21706
rect 219 21658 1619 21664
rect 1660 21660 1706 21672
rect 219 21624 231 21658
rect 1607 21624 1619 21658
rect 132 21610 178 21622
rect 219 21618 1619 21624
rect 132 21576 138 21610
rect 172 21576 178 21610
rect 132 21564 178 21576
rect 219 21562 1619 21568
rect 219 21528 231 21562
rect 1607 21528 1619 21562
rect 219 21522 1619 21528
rect 1660 21514 1706 21526
rect 1660 21480 1666 21514
rect 1700 21480 1706 21514
rect 219 21466 1619 21472
rect 1660 21468 1706 21480
rect 219 21432 231 21466
rect 1607 21432 1619 21466
rect 132 21418 178 21430
rect 219 21426 1619 21432
rect 132 21384 138 21418
rect 172 21384 178 21418
rect 132 21372 178 21384
rect 219 21370 1619 21376
rect 219 21336 231 21370
rect 1607 21336 1619 21370
rect 219 21330 1619 21336
rect 1660 21322 1706 21334
rect 1660 21288 1666 21322
rect 1700 21288 1706 21322
rect 219 21274 1619 21280
rect 1660 21276 1706 21288
rect 219 21240 231 21274
rect 1607 21240 1619 21274
rect 132 21226 178 21238
rect 219 21234 1619 21240
rect 132 21192 138 21226
rect 172 21192 178 21226
rect 132 21180 178 21192
rect 219 21178 1619 21184
rect 219 21144 231 21178
rect 1607 21144 1619 21178
rect 219 21138 1619 21144
rect 1660 21130 1706 21142
rect 1660 21096 1666 21130
rect 1700 21096 1706 21130
rect 219 21082 1619 21088
rect 1660 21084 1706 21096
rect 219 21048 231 21082
rect 1607 21048 1619 21082
rect 132 21034 178 21046
rect 219 21042 1619 21048
rect 132 21000 138 21034
rect 172 21000 178 21034
rect 132 20988 178 21000
rect 219 20986 1619 20992
rect 219 20952 231 20986
rect 1607 20952 1619 20986
rect 219 20946 1619 20952
rect 1660 20938 1706 20950
rect 1660 20904 1666 20938
rect 1700 20904 1706 20938
rect 219 20890 1619 20896
rect 1660 20892 1706 20904
rect 219 20856 231 20890
rect 1607 20856 1619 20890
rect 132 20842 178 20854
rect 219 20850 1619 20856
rect 132 20808 138 20842
rect 172 20808 178 20842
rect 132 20796 178 20808
rect 219 20794 1619 20800
rect 219 20760 231 20794
rect 1607 20760 1619 20794
rect 219 20754 1619 20760
rect 1660 20746 1706 20758
rect 1660 20712 1666 20746
rect 1700 20712 1706 20746
rect 219 20698 1619 20704
rect 1660 20700 1706 20712
rect 219 20664 231 20698
rect 1607 20664 1619 20698
rect 132 20650 178 20662
rect 219 20658 1619 20664
rect 132 20616 138 20650
rect 172 20616 178 20650
rect 132 20604 178 20616
rect 219 20602 1619 20608
rect 219 20568 231 20602
rect 1607 20568 1619 20602
rect 219 20562 1619 20568
rect 1660 20554 1706 20566
rect 1660 20520 1666 20554
rect 1700 20520 1706 20554
rect 219 20506 1619 20512
rect 1660 20508 1706 20520
rect 219 20472 231 20506
rect 1607 20472 1619 20506
rect 132 20458 178 20470
rect 219 20466 1619 20472
rect 132 20424 138 20458
rect 172 20424 178 20458
rect 132 20412 178 20424
rect 219 20410 1619 20416
rect 219 20376 231 20410
rect 1607 20376 1619 20410
rect 219 20370 1619 20376
rect 1660 20362 1706 20374
rect 1660 20328 1666 20362
rect 1700 20328 1706 20362
rect 219 20314 1619 20320
rect 1660 20316 1706 20328
rect 219 20280 231 20314
rect 1607 20280 1619 20314
rect 132 20266 178 20278
rect 219 20274 1619 20280
rect 132 20232 138 20266
rect 172 20232 178 20266
rect 132 20220 178 20232
rect 219 20218 1619 20224
rect 219 20184 231 20218
rect 1607 20184 1619 20218
rect 219 20178 1619 20184
rect 1660 20170 1706 20182
rect 1660 20136 1666 20170
rect 1700 20136 1706 20170
rect 219 20122 1619 20128
rect 1660 20124 1706 20136
rect 219 20088 231 20122
rect 1607 20088 1619 20122
rect 132 20074 178 20086
rect 219 20082 1619 20088
rect 132 20040 138 20074
rect 172 20040 178 20074
rect 132 20028 178 20040
rect 219 20026 1619 20032
rect 219 19992 231 20026
rect 1607 19992 1619 20026
rect 219 19986 1619 19992
rect 1660 19978 1706 19990
rect 1660 19944 1666 19978
rect 1700 19944 1706 19978
rect 219 19930 1619 19936
rect 1660 19932 1706 19944
rect 219 19896 231 19930
rect 1607 19896 1619 19930
rect 132 19882 178 19894
rect 219 19890 1619 19896
rect 132 19848 138 19882
rect 172 19848 178 19882
rect 132 19836 178 19848
rect 219 19834 1619 19840
rect 219 19800 231 19834
rect 1607 19800 1619 19834
rect 219 19794 1619 19800
rect 1660 19786 1706 19798
rect 1660 19752 1666 19786
rect 1700 19752 1706 19786
rect 219 19738 1619 19744
rect 1660 19740 1706 19752
rect 219 19704 231 19738
rect 1607 19704 1619 19738
rect 132 19690 178 19702
rect 219 19698 1619 19704
rect 132 19656 138 19690
rect 172 19656 178 19690
rect 132 19644 178 19656
rect 219 19642 1619 19648
rect 219 19608 231 19642
rect 1607 19608 1619 19642
rect 219 19602 1619 19608
rect 1660 19594 1706 19606
rect 1660 19560 1666 19594
rect 1700 19560 1706 19594
rect 219 19546 1619 19552
rect 1660 19548 1706 19560
rect 219 19512 231 19546
rect 1607 19512 1619 19546
rect 132 19498 178 19510
rect 219 19506 1619 19512
rect 132 19464 138 19498
rect 172 19464 178 19498
rect 132 19452 178 19464
rect 219 19450 1619 19456
rect 219 19416 231 19450
rect 1607 19416 1619 19450
rect 219 19410 1619 19416
rect 1660 19402 1706 19414
rect 1660 19368 1666 19402
rect 1700 19368 1706 19402
rect 219 19354 1619 19360
rect 1660 19356 1706 19368
rect 219 19320 231 19354
rect 1607 19320 1619 19354
rect 132 19306 178 19318
rect 219 19314 1619 19320
rect 132 19272 138 19306
rect 172 19272 178 19306
rect 132 19260 178 19272
rect 219 19258 1619 19264
rect 219 19224 231 19258
rect 1607 19224 1619 19258
rect 219 19218 1619 19224
rect 1660 19210 1706 19222
rect 1660 19176 1666 19210
rect 1700 19176 1706 19210
rect 219 19162 1619 19168
rect 1660 19164 1706 19176
rect 219 19128 231 19162
rect 1607 19128 1619 19162
rect 132 19114 178 19126
rect 219 19122 1619 19128
rect 132 19080 138 19114
rect 172 19080 178 19114
rect 132 19068 178 19080
rect 219 19066 1619 19072
rect 219 19032 231 19066
rect 1607 19032 1619 19066
rect 219 19026 1619 19032
rect 1660 19018 1706 19030
rect 1660 18984 1666 19018
rect 1700 18984 1706 19018
rect 219 18970 1619 18976
rect 1660 18972 1706 18984
rect 219 18936 231 18970
rect 1607 18936 1619 18970
rect 132 18922 178 18934
rect 219 18930 1619 18936
rect 132 18888 138 18922
rect 172 18888 178 18922
rect 132 18876 178 18888
rect 219 18874 1619 18880
rect 219 18840 231 18874
rect 1607 18840 1619 18874
rect 219 18834 1619 18840
rect 1660 18826 1706 18838
rect 1660 18792 1666 18826
rect 1700 18792 1706 18826
rect 219 18778 1619 18784
rect 1660 18780 1706 18792
rect 219 18744 231 18778
rect 1607 18744 1619 18778
rect 132 18730 178 18742
rect 219 18738 1619 18744
rect 132 18696 138 18730
rect 172 18696 178 18730
rect 132 18684 178 18696
rect 219 18682 1619 18688
rect 219 18648 231 18682
rect 1607 18648 1619 18682
rect 219 18642 1619 18648
rect 1660 18634 1706 18646
rect 1660 18600 1666 18634
rect 1700 18600 1706 18634
rect 219 18586 1619 18592
rect 1660 18588 1706 18600
rect 219 18552 231 18586
rect 1607 18552 1619 18586
rect 132 18538 178 18550
rect 219 18546 1619 18552
rect 132 18504 138 18538
rect 172 18504 178 18538
rect 132 18492 178 18504
rect 219 18490 1619 18496
rect 219 18456 231 18490
rect 1607 18456 1619 18490
rect 219 18450 1619 18456
rect 1660 18442 1706 18454
rect 1660 18408 1666 18442
rect 1700 18408 1706 18442
rect 219 18394 1619 18400
rect 1660 18396 1706 18408
rect 219 18360 231 18394
rect 1607 18360 1619 18394
rect 132 18346 178 18358
rect 219 18354 1619 18360
rect 132 18312 138 18346
rect 172 18312 178 18346
rect 132 18300 178 18312
rect 219 18298 1619 18304
rect 219 18264 231 18298
rect 1607 18264 1619 18298
rect 219 18258 1619 18264
rect 1660 18250 1706 18262
rect 1660 18216 1666 18250
rect 1700 18216 1706 18250
rect 219 18202 1619 18208
rect 1660 18204 1706 18216
rect 219 18168 231 18202
rect 1607 18168 1619 18202
rect 132 18154 178 18166
rect 219 18162 1619 18168
rect 132 18120 138 18154
rect 172 18120 178 18154
rect 132 18108 178 18120
rect 219 18106 1619 18112
rect 219 18072 231 18106
rect 1607 18072 1619 18106
rect 219 18066 1619 18072
rect 1660 18058 1706 18070
rect 1660 18024 1666 18058
rect 1700 18024 1706 18058
rect 219 18010 1619 18016
rect 1660 18012 1706 18024
rect 219 17976 231 18010
rect 1607 17976 1619 18010
rect 132 17962 178 17974
rect 219 17970 1619 17976
rect 132 17928 138 17962
rect 172 17928 178 17962
rect 132 17916 178 17928
rect 219 17914 1619 17920
rect 219 17880 231 17914
rect 1607 17880 1619 17914
rect 219 17874 1619 17880
rect 1660 17866 1706 17878
rect 1660 17832 1666 17866
rect 1700 17832 1706 17866
rect 219 17818 1619 17824
rect 1660 17820 1706 17832
rect 219 17784 231 17818
rect 1607 17784 1619 17818
rect 132 17770 178 17782
rect 219 17778 1619 17784
rect 132 17736 138 17770
rect 172 17736 178 17770
rect 132 17724 178 17736
rect 219 17722 1619 17728
rect 219 17688 231 17722
rect 1607 17688 1619 17722
rect 219 17682 1619 17688
rect 1660 17674 1706 17686
rect 1660 17640 1666 17674
rect 1700 17640 1706 17674
rect 219 17626 1619 17632
rect 1660 17628 1706 17640
rect 219 17592 231 17626
rect 1607 17592 1619 17626
rect 132 17578 178 17590
rect 219 17586 1619 17592
rect 132 17544 138 17578
rect 172 17544 178 17578
rect 132 17532 178 17544
rect 219 17530 1619 17536
rect 219 17496 231 17530
rect 1607 17496 1619 17530
rect 219 17490 1619 17496
rect 1660 17482 1706 17494
rect 1660 17448 1666 17482
rect 1700 17448 1706 17482
rect 219 17434 1619 17440
rect 1660 17436 1706 17448
rect 219 17400 231 17434
rect 1607 17400 1619 17434
rect 132 17386 178 17398
rect 219 17394 1619 17400
rect 132 17352 138 17386
rect 172 17352 178 17386
rect 132 17340 178 17352
rect 219 17338 1619 17344
rect 219 17304 231 17338
rect 1607 17304 1619 17338
rect 219 17298 1619 17304
rect 1660 17290 1706 17302
rect 1660 17256 1666 17290
rect 1700 17256 1706 17290
rect 219 17242 1619 17248
rect 1660 17244 1706 17256
rect 219 17208 231 17242
rect 1607 17208 1619 17242
rect 132 17194 178 17206
rect 219 17202 1619 17208
rect 132 17160 138 17194
rect 172 17160 178 17194
rect 132 17148 178 17160
rect 219 17146 1619 17152
rect 219 17112 231 17146
rect 1607 17112 1619 17146
rect 219 17106 1619 17112
rect 1660 17098 1706 17110
rect 1660 17064 1666 17098
rect 1700 17064 1706 17098
rect 219 17050 1619 17056
rect 1660 17052 1706 17064
rect 219 17016 231 17050
rect 1607 17016 1619 17050
rect 132 17002 178 17014
rect 219 17010 1619 17016
rect 132 16968 138 17002
rect 172 16968 178 17002
rect 132 16956 178 16968
rect 219 16954 1619 16960
rect 219 16920 231 16954
rect 1607 16920 1619 16954
rect 219 16914 1619 16920
rect 1660 16906 1706 16918
rect 1660 16872 1666 16906
rect 1700 16872 1706 16906
rect 219 16858 1619 16864
rect 1660 16860 1706 16872
rect 219 16824 231 16858
rect 1607 16824 1619 16858
rect 132 16810 178 16822
rect 219 16818 1619 16824
rect 132 16776 138 16810
rect 172 16776 178 16810
rect 132 16764 178 16776
rect 219 16762 1619 16768
rect 219 16728 231 16762
rect 1607 16728 1619 16762
rect 219 16722 1619 16728
rect 1660 16714 1706 16726
rect 1660 16680 1666 16714
rect 1700 16680 1706 16714
rect 219 16666 1619 16672
rect 1660 16668 1706 16680
rect 219 16632 231 16666
rect 1607 16632 1619 16666
rect 132 16618 178 16630
rect 219 16626 1619 16632
rect 132 16584 138 16618
rect 172 16584 178 16618
rect 132 16572 178 16584
rect 219 16570 1619 16576
rect 219 16536 231 16570
rect 1607 16536 1619 16570
rect 219 16530 1619 16536
rect 1660 16522 1706 16534
rect 1660 16488 1666 16522
rect 1700 16488 1706 16522
rect 219 16474 1619 16480
rect 1660 16476 1706 16488
rect 219 16440 231 16474
rect 1607 16440 1619 16474
rect 132 16426 178 16438
rect 219 16434 1619 16440
rect 132 16392 138 16426
rect 172 16392 178 16426
rect 132 16380 178 16392
rect 219 16378 1619 16384
rect 219 16344 231 16378
rect 1607 16344 1619 16378
rect 219 16338 1619 16344
rect 1660 16330 1706 16342
rect 1660 16296 1666 16330
rect 1700 16296 1706 16330
rect 219 16282 1619 16288
rect 1660 16284 1706 16296
rect 219 16248 231 16282
rect 1607 16248 1619 16282
rect 132 16234 178 16246
rect 219 16242 1619 16248
rect 132 16200 138 16234
rect 172 16200 178 16234
rect 132 16188 178 16200
rect 219 16186 1619 16192
rect 219 16152 231 16186
rect 1607 16152 1619 16186
rect 219 16146 1619 16152
rect 1660 16138 1706 16150
rect 1660 16104 1666 16138
rect 1700 16104 1706 16138
rect 219 16090 1619 16096
rect 1660 16092 1706 16104
rect 219 16056 231 16090
rect 1607 16056 1619 16090
rect 132 16042 178 16054
rect 219 16050 1619 16056
rect 132 16008 138 16042
rect 172 16008 178 16042
rect 132 15996 178 16008
rect 219 15994 1619 16000
rect 219 15960 231 15994
rect 1607 15960 1619 15994
rect 219 15954 1619 15960
rect 1660 15946 1706 15958
rect 1660 15912 1666 15946
rect 1700 15912 1706 15946
rect 219 15898 1619 15904
rect 1660 15900 1706 15912
rect 219 15864 231 15898
rect 1607 15864 1619 15898
rect 132 15850 178 15862
rect 219 15858 1619 15864
rect 132 15816 138 15850
rect 172 15816 178 15850
rect 132 15804 178 15816
rect 219 15802 1619 15808
rect 219 15768 231 15802
rect 1607 15768 1619 15802
rect 219 15762 1619 15768
rect 1660 15754 1706 15766
rect 1660 15720 1666 15754
rect 1700 15720 1706 15754
rect 219 15706 1619 15712
rect 1660 15708 1706 15720
rect 219 15672 231 15706
rect 1607 15672 1619 15706
rect 132 15658 178 15670
rect 219 15666 1619 15672
rect 132 15624 138 15658
rect 172 15624 178 15658
rect 132 15612 178 15624
rect 219 15610 1619 15616
rect 219 15576 231 15610
rect 1607 15576 1619 15610
rect 219 15570 1619 15576
rect 1660 15562 1706 15574
rect 1660 15528 1666 15562
rect 1700 15528 1706 15562
rect 219 15514 1619 15520
rect 1660 15516 1706 15528
rect 219 15480 231 15514
rect 1607 15480 1619 15514
rect 132 15466 178 15478
rect 219 15474 1619 15480
rect 132 15432 138 15466
rect 172 15432 178 15466
rect 132 15420 178 15432
rect 219 15418 1619 15424
rect 219 15384 231 15418
rect 1607 15384 1619 15418
rect 219 15378 1619 15384
rect 1660 15370 1706 15382
rect 1660 15336 1666 15370
rect 1700 15336 1706 15370
rect 219 15322 1619 15328
rect 1660 15324 1706 15336
rect 219 15288 231 15322
rect 1607 15288 1619 15322
rect 132 15274 178 15286
rect 219 15282 1619 15288
rect 132 15240 138 15274
rect 172 15240 178 15274
rect 132 15228 178 15240
rect 219 15226 1619 15232
rect 219 15192 231 15226
rect 1607 15192 1619 15226
rect 219 15186 1619 15192
rect 1660 15178 1706 15190
rect 1660 15144 1666 15178
rect 1700 15144 1706 15178
rect 219 15130 1619 15136
rect 1660 15132 1706 15144
rect 219 15096 231 15130
rect 1607 15096 1619 15130
rect 132 15082 178 15094
rect 219 15090 1619 15096
rect 132 15048 138 15082
rect 172 15048 178 15082
rect 132 15036 178 15048
rect 219 15034 1619 15040
rect 219 15000 231 15034
rect 1607 15000 1619 15034
rect 219 14994 1619 15000
rect 1660 14986 1706 14998
rect 1660 14952 1666 14986
rect 1700 14952 1706 14986
rect 219 14938 1619 14944
rect 1660 14940 1706 14952
rect 219 14904 231 14938
rect 1607 14904 1619 14938
rect 132 14890 178 14902
rect 219 14898 1619 14904
rect 132 14856 138 14890
rect 172 14856 178 14890
rect 132 14844 178 14856
rect 219 14842 1619 14848
rect 219 14808 231 14842
rect 1607 14808 1619 14842
rect 219 14802 1619 14808
rect 1660 14794 1706 14806
rect 1660 14760 1666 14794
rect 1700 14760 1706 14794
rect 219 14746 1619 14752
rect 1660 14748 1706 14760
rect 219 14712 231 14746
rect 1607 14712 1619 14746
rect 132 14698 178 14710
rect 219 14706 1619 14712
rect 132 14664 138 14698
rect 172 14664 178 14698
rect 132 14652 178 14664
rect 219 14650 1619 14656
rect 219 14616 231 14650
rect 1607 14616 1619 14650
rect 219 14610 1619 14616
rect 1660 14602 1706 14614
rect 1660 14568 1666 14602
rect 1700 14568 1706 14602
rect 219 14554 1619 14560
rect 1660 14556 1706 14568
rect 219 14520 231 14554
rect 1607 14520 1619 14554
rect 132 14506 178 14518
rect 219 14514 1619 14520
rect 132 14472 138 14506
rect 172 14472 178 14506
rect 132 14460 178 14472
rect 219 14458 1619 14464
rect 219 14424 231 14458
rect 1607 14424 1619 14458
rect 219 14418 1619 14424
rect 1660 14410 1706 14422
rect 1660 14376 1666 14410
rect 1700 14376 1706 14410
rect 219 14362 1619 14368
rect 1660 14364 1706 14376
rect 219 14328 231 14362
rect 1607 14328 1619 14362
rect 132 14314 178 14326
rect 219 14322 1619 14328
rect 132 14280 138 14314
rect 172 14280 178 14314
rect 132 14268 178 14280
rect 219 14266 1619 14272
rect 219 14232 231 14266
rect 1607 14232 1619 14266
rect 219 14226 1619 14232
rect 1660 14218 1706 14230
rect 1660 14184 1666 14218
rect 1700 14184 1706 14218
rect 219 14170 1619 14176
rect 1660 14172 1706 14184
rect 219 14136 231 14170
rect 1607 14136 1619 14170
rect 132 14122 178 14134
rect 219 14130 1619 14136
rect 132 14088 138 14122
rect 172 14088 178 14122
rect 132 14076 178 14088
rect 219 14074 1619 14080
rect 219 14040 231 14074
rect 1607 14040 1619 14074
rect 219 14034 1619 14040
rect 1660 14026 1706 14038
rect 1660 13992 1666 14026
rect 1700 13992 1706 14026
rect 219 13978 1619 13984
rect 1660 13980 1706 13992
rect 219 13944 231 13978
rect 1607 13944 1619 13978
rect 132 13930 178 13942
rect 219 13938 1619 13944
rect 132 13896 138 13930
rect 172 13896 178 13930
rect 132 13884 178 13896
rect 219 13882 1619 13888
rect 219 13848 231 13882
rect 1607 13848 1619 13882
rect 219 13842 1619 13848
rect 1660 13834 1706 13846
rect 1660 13800 1666 13834
rect 1700 13800 1706 13834
rect 219 13786 1619 13792
rect 1660 13788 1706 13800
rect 219 13752 231 13786
rect 1607 13752 1619 13786
rect 132 13738 178 13750
rect 219 13746 1619 13752
rect 132 13704 138 13738
rect 172 13704 178 13738
rect 132 13692 178 13704
rect 219 13690 1619 13696
rect 219 13656 231 13690
rect 1607 13656 1619 13690
rect 219 13650 1619 13656
rect 1660 13642 1706 13654
rect 1660 13608 1666 13642
rect 1700 13608 1706 13642
rect 219 13594 1619 13600
rect 1660 13596 1706 13608
rect 219 13560 231 13594
rect 1607 13560 1619 13594
rect 132 13546 178 13558
rect 219 13554 1619 13560
rect 132 13512 138 13546
rect 172 13512 178 13546
rect 132 13500 178 13512
rect 219 13498 1619 13504
rect 219 13464 231 13498
rect 1607 13464 1619 13498
rect 219 13458 1619 13464
rect 1660 13450 1706 13462
rect 1660 13416 1666 13450
rect 1700 13416 1706 13450
rect 219 13402 1619 13408
rect 1660 13404 1706 13416
rect 219 13368 231 13402
rect 1607 13368 1619 13402
rect 132 13354 178 13366
rect 219 13362 1619 13368
rect 132 13320 138 13354
rect 172 13320 178 13354
rect 132 13308 178 13320
rect 219 13306 1619 13312
rect 219 13272 231 13306
rect 1607 13272 1619 13306
rect 219 13266 1619 13272
rect 1660 13258 1706 13270
rect 1660 13224 1666 13258
rect 1700 13224 1706 13258
rect 219 13210 1619 13216
rect 1660 13212 1706 13224
rect 219 13176 231 13210
rect 1607 13176 1619 13210
rect 132 13162 178 13174
rect 219 13170 1619 13176
rect 132 13128 138 13162
rect 172 13128 178 13162
rect 132 13116 178 13128
rect 219 13114 1619 13120
rect 219 13080 231 13114
rect 1607 13080 1619 13114
rect 219 13074 1619 13080
rect 1660 13066 1706 13078
rect 1660 13032 1666 13066
rect 1700 13032 1706 13066
rect 219 13018 1619 13024
rect 1660 13020 1706 13032
rect 219 12984 231 13018
rect 1607 12984 1619 13018
rect 132 12970 178 12982
rect 219 12978 1619 12984
rect 132 12936 138 12970
rect 172 12936 178 12970
rect 132 12924 178 12936
rect 219 12922 1619 12928
rect 219 12888 231 12922
rect 1607 12888 1619 12922
rect 219 12882 1619 12888
rect 1660 12874 1706 12886
rect 1660 12840 1666 12874
rect 1700 12840 1706 12874
rect 219 12826 1619 12832
rect 1660 12828 1706 12840
rect 219 12792 231 12826
rect 1607 12792 1619 12826
rect 132 12778 178 12790
rect 219 12786 1619 12792
rect 132 12744 138 12778
rect 172 12744 178 12778
rect 132 12732 178 12744
rect 219 12730 1619 12736
rect 219 12696 231 12730
rect 1607 12696 1619 12730
rect 219 12690 1619 12696
rect 1660 12682 1706 12694
rect 1660 12648 1666 12682
rect 1700 12648 1706 12682
rect 219 12634 1619 12640
rect 1660 12636 1706 12648
rect 219 12600 231 12634
rect 1607 12600 1619 12634
rect 132 12586 178 12598
rect 219 12594 1619 12600
rect 132 12552 138 12586
rect 172 12552 178 12586
rect 132 12540 178 12552
rect 219 12538 1619 12544
rect 219 12504 231 12538
rect 1607 12504 1619 12538
rect 219 12498 1619 12504
rect 1660 12490 1706 12502
rect 1660 12456 1666 12490
rect 1700 12456 1706 12490
rect 219 12442 1619 12448
rect 1660 12444 1706 12456
rect 219 12408 231 12442
rect 1607 12408 1619 12442
rect 132 12394 178 12406
rect 219 12402 1619 12408
rect 132 12360 138 12394
rect 172 12360 178 12394
rect 132 12348 178 12360
rect 219 12346 1619 12352
rect 219 12312 231 12346
rect 1607 12312 1619 12346
rect 219 12306 1619 12312
rect 1660 12298 1706 12310
rect 1660 12264 1666 12298
rect 1700 12264 1706 12298
rect 219 12250 1619 12256
rect 1660 12252 1706 12264
rect 219 12216 231 12250
rect 1607 12216 1619 12250
rect 132 12202 178 12214
rect 219 12210 1619 12216
rect 132 12168 138 12202
rect 172 12168 178 12202
rect 132 12156 178 12168
rect 219 12154 1619 12160
rect 219 12120 231 12154
rect 1607 12120 1619 12154
rect 219 12114 1619 12120
rect 1660 12106 1706 12118
rect 1660 12072 1666 12106
rect 1700 12072 1706 12106
rect 219 12058 1619 12064
rect 1660 12060 1706 12072
rect 219 12024 231 12058
rect 1607 12024 1619 12058
rect 132 12010 178 12022
rect 219 12018 1619 12024
rect 132 11976 138 12010
rect 172 11976 178 12010
rect 132 11964 178 11976
rect 219 11962 1619 11968
rect 219 11928 231 11962
rect 1607 11928 1619 11962
rect 219 11922 1619 11928
rect 1660 11914 1706 11926
rect 1660 11880 1666 11914
rect 1700 11880 1706 11914
rect 219 11866 1619 11872
rect 1660 11868 1706 11880
rect 219 11832 231 11866
rect 1607 11832 1619 11866
rect 132 11818 178 11830
rect 219 11826 1619 11832
rect 132 11784 138 11818
rect 172 11784 178 11818
rect 132 11772 178 11784
rect 219 11770 1619 11776
rect 219 11736 231 11770
rect 1607 11736 1619 11770
rect 219 11730 1619 11736
rect 1660 11722 1706 11734
rect 1660 11688 1666 11722
rect 1700 11688 1706 11722
rect 219 11674 1619 11680
rect 1660 11676 1706 11688
rect 219 11640 231 11674
rect 1607 11640 1619 11674
rect 132 11626 178 11638
rect 219 11634 1619 11640
rect 132 11592 138 11626
rect 172 11592 178 11626
rect 132 11580 178 11592
rect 219 11578 1619 11584
rect 219 11544 231 11578
rect 1607 11544 1619 11578
rect 219 11538 1619 11544
rect 1660 11530 1706 11542
rect 1660 11496 1666 11530
rect 1700 11496 1706 11530
rect 219 11482 1619 11488
rect 1660 11484 1706 11496
rect 219 11448 231 11482
rect 1607 11448 1619 11482
rect 132 11434 178 11446
rect 219 11442 1619 11448
rect 132 11400 138 11434
rect 172 11400 178 11434
rect 132 11388 178 11400
rect 219 11386 1619 11392
rect 219 11352 231 11386
rect 1607 11352 1619 11386
rect 219 11346 1619 11352
rect 1660 11338 1706 11350
rect 1660 11304 1666 11338
rect 1700 11304 1706 11338
rect 219 11290 1619 11296
rect 1660 11292 1706 11304
rect 219 11256 231 11290
rect 1607 11256 1619 11290
rect 132 11242 178 11254
rect 219 11250 1619 11256
rect 132 11208 138 11242
rect 172 11208 178 11242
rect 132 11196 178 11208
rect 219 11194 1619 11200
rect 219 11160 231 11194
rect 1607 11160 1619 11194
rect 219 11154 1619 11160
rect 1660 11146 1706 11158
rect 1660 11112 1666 11146
rect 1700 11112 1706 11146
rect 219 11098 1619 11104
rect 1660 11100 1706 11112
rect 219 11064 231 11098
rect 1607 11064 1619 11098
rect 132 11050 178 11062
rect 219 11058 1619 11064
rect 132 11016 138 11050
rect 172 11016 178 11050
rect 132 11004 178 11016
rect 219 11002 1619 11008
rect 219 10968 231 11002
rect 1607 10968 1619 11002
rect 219 10962 1619 10968
rect 1660 10954 1706 10966
rect 1660 10920 1666 10954
rect 1700 10920 1706 10954
rect 219 10906 1619 10912
rect 1660 10908 1706 10920
rect 219 10872 231 10906
rect 1607 10872 1619 10906
rect 132 10858 178 10870
rect 219 10866 1619 10872
rect 132 10824 138 10858
rect 172 10824 178 10858
rect 132 10812 178 10824
rect 219 10810 1619 10816
rect 219 10776 231 10810
rect 1607 10776 1619 10810
rect 219 10770 1619 10776
rect 1660 10762 1706 10774
rect 1660 10728 1666 10762
rect 1700 10728 1706 10762
rect 219 10714 1619 10720
rect 1660 10716 1706 10728
rect 219 10680 231 10714
rect 1607 10680 1619 10714
rect 132 10666 178 10678
rect 219 10674 1619 10680
rect 132 10632 138 10666
rect 172 10632 178 10666
rect 132 10620 178 10632
rect 219 10618 1619 10624
rect 219 10584 231 10618
rect 1607 10584 1619 10618
rect 219 10578 1619 10584
rect 1660 10570 1706 10582
rect 1660 10536 1666 10570
rect 1700 10536 1706 10570
rect 219 10522 1619 10528
rect 1660 10524 1706 10536
rect 219 10488 231 10522
rect 1607 10488 1619 10522
rect 132 10474 178 10486
rect 219 10482 1619 10488
rect 132 10440 138 10474
rect 172 10440 178 10474
rect 132 10428 178 10440
rect 219 10426 1619 10432
rect 219 10392 231 10426
rect 1607 10392 1619 10426
rect 219 10386 1619 10392
rect 1660 10378 1706 10390
rect 1660 10344 1666 10378
rect 1700 10344 1706 10378
rect 219 10330 1619 10336
rect 1660 10332 1706 10344
rect 219 10296 231 10330
rect 1607 10296 1619 10330
rect 132 10282 178 10294
rect 219 10290 1619 10296
rect 132 10248 138 10282
rect 172 10248 178 10282
rect 132 10236 178 10248
rect 219 10234 1619 10240
rect 219 10200 231 10234
rect 1607 10200 1619 10234
rect 219 10194 1619 10200
rect 1660 10186 1706 10198
rect 1660 10152 1666 10186
rect 1700 10152 1706 10186
rect 219 10138 1619 10144
rect 1660 10140 1706 10152
rect 219 10104 231 10138
rect 1607 10104 1619 10138
rect 132 10090 178 10102
rect 219 10098 1619 10104
rect 132 10056 138 10090
rect 172 10056 178 10090
rect 132 10044 178 10056
rect 219 10042 1619 10048
rect 219 10008 231 10042
rect 1607 10008 1619 10042
rect 219 10002 1619 10008
rect 1660 9994 1706 10006
rect 1660 9960 1666 9994
rect 1700 9960 1706 9994
rect 219 9946 1619 9952
rect 1660 9948 1706 9960
rect 219 9912 231 9946
rect 1607 9912 1619 9946
rect 132 9898 178 9910
rect 219 9906 1619 9912
rect 132 9864 138 9898
rect 172 9864 178 9898
rect 132 9852 178 9864
rect 219 9850 1619 9856
rect 219 9816 231 9850
rect 1607 9816 1619 9850
rect 219 9810 1619 9816
rect 1660 9802 1706 9814
rect 1660 9768 1666 9802
rect 1700 9768 1706 9802
rect 219 9754 1619 9760
rect 1660 9756 1706 9768
rect 219 9720 231 9754
rect 1607 9720 1619 9754
rect 132 9706 178 9718
rect 219 9714 1619 9720
rect 132 9672 138 9706
rect 172 9672 178 9706
rect 132 9660 178 9672
rect 219 9658 1619 9664
rect 219 9624 231 9658
rect 1607 9624 1619 9658
rect 219 9618 1619 9624
rect 1660 9610 1706 9622
rect 1660 9576 1666 9610
rect 1700 9576 1706 9610
rect 219 9562 1619 9568
rect 1660 9564 1706 9576
rect 219 9528 231 9562
rect 1607 9528 1619 9562
rect 132 9514 178 9526
rect 219 9522 1619 9528
rect 132 9480 138 9514
rect 172 9480 178 9514
rect 132 9468 178 9480
rect 219 9466 1619 9472
rect 219 9432 231 9466
rect 1607 9432 1619 9466
rect 219 9426 1619 9432
rect 1660 9418 1706 9430
rect 1660 9384 1666 9418
rect 1700 9384 1706 9418
rect 219 9370 1619 9376
rect 1660 9372 1706 9384
rect 219 9336 231 9370
rect 1607 9336 1619 9370
rect 132 9322 178 9334
rect 219 9330 1619 9336
rect 132 9288 138 9322
rect 172 9288 178 9322
rect 132 9276 178 9288
rect 219 9274 1619 9280
rect 219 9240 231 9274
rect 1607 9240 1619 9274
rect 219 9234 1619 9240
rect 1660 9226 1706 9238
rect 1660 9192 1666 9226
rect 1700 9192 1706 9226
rect 219 9178 1619 9184
rect 1660 9180 1706 9192
rect 219 9144 231 9178
rect 1607 9144 1619 9178
rect 132 9130 178 9142
rect 219 9138 1619 9144
rect 132 9096 138 9130
rect 172 9096 178 9130
rect 132 9084 178 9096
rect 219 9082 1619 9088
rect 219 9048 231 9082
rect 1607 9048 1619 9082
rect 219 9042 1619 9048
rect 1660 9034 1706 9046
rect 1660 9000 1666 9034
rect 1700 9000 1706 9034
rect 219 8986 1619 8992
rect 1660 8988 1706 9000
rect 219 8952 231 8986
rect 1607 8952 1619 8986
rect 132 8938 178 8950
rect 219 8946 1619 8952
rect 132 8904 138 8938
rect 172 8904 178 8938
rect 132 8892 178 8904
rect 219 8890 1619 8896
rect 219 8856 231 8890
rect 1607 8856 1619 8890
rect 219 8850 1619 8856
rect 1660 8842 1706 8854
rect 1660 8808 1666 8842
rect 1700 8808 1706 8842
rect 219 8794 1619 8800
rect 1660 8796 1706 8808
rect 219 8760 231 8794
rect 1607 8760 1619 8794
rect 132 8746 178 8758
rect 219 8754 1619 8760
rect 132 8712 138 8746
rect 172 8712 178 8746
rect 132 8700 178 8712
rect 219 8698 1619 8704
rect 219 8664 231 8698
rect 1607 8664 1619 8698
rect 219 8658 1619 8664
rect 1660 8650 1706 8662
rect 1660 8616 1666 8650
rect 1700 8616 1706 8650
rect 219 8602 1619 8608
rect 1660 8604 1706 8616
rect 219 8568 231 8602
rect 1607 8568 1619 8602
rect 132 8554 178 8566
rect 219 8562 1619 8568
rect 132 8520 138 8554
rect 172 8520 178 8554
rect 132 8508 178 8520
rect 219 8506 1619 8512
rect 219 8472 231 8506
rect 1607 8472 1619 8506
rect 219 8466 1619 8472
rect 1660 8458 1706 8470
rect 1660 8424 1666 8458
rect 1700 8424 1706 8458
rect 219 8410 1619 8416
rect 1660 8412 1706 8424
rect 219 8376 231 8410
rect 1607 8376 1619 8410
rect 132 8362 178 8374
rect 219 8370 1619 8376
rect 132 8328 138 8362
rect 172 8328 178 8362
rect 132 8316 178 8328
rect 219 8314 1619 8320
rect 219 8280 231 8314
rect 1607 8280 1619 8314
rect 219 8274 1619 8280
rect 1660 8266 1706 8278
rect 1660 8232 1666 8266
rect 1700 8232 1706 8266
rect 219 8218 1619 8224
rect 1660 8220 1706 8232
rect 219 8184 231 8218
rect 1607 8184 1619 8218
rect 132 8170 178 8182
rect 219 8178 1619 8184
rect 132 8136 138 8170
rect 172 8136 178 8170
rect 132 8124 178 8136
rect 219 8122 1619 8128
rect 219 8088 231 8122
rect 1607 8088 1619 8122
rect 219 8082 1619 8088
rect 1660 8074 1706 8086
rect 1660 8040 1666 8074
rect 1700 8040 1706 8074
rect 219 8026 1619 8032
rect 1660 8028 1706 8040
rect 219 7992 231 8026
rect 1607 7992 1619 8026
rect 132 7978 178 7990
rect 219 7986 1619 7992
rect 132 7944 138 7978
rect 172 7944 178 7978
rect 132 7932 178 7944
rect 219 7930 1619 7936
rect 219 7896 231 7930
rect 1607 7896 1619 7930
rect 219 7890 1619 7896
rect 1660 7882 1706 7894
rect 1660 7848 1666 7882
rect 1700 7848 1706 7882
rect 219 7834 1619 7840
rect 1660 7836 1706 7848
rect 219 7800 231 7834
rect 1607 7800 1619 7834
rect 132 7786 178 7798
rect 219 7794 1619 7800
rect 132 7752 138 7786
rect 172 7752 178 7786
rect 132 7740 178 7752
rect 219 7738 1619 7744
rect 219 7704 231 7738
rect 1607 7704 1619 7738
rect 219 7698 1619 7704
rect 1660 7690 1706 7702
rect 1660 7656 1666 7690
rect 1700 7656 1706 7690
rect 219 7642 1619 7648
rect 1660 7644 1706 7656
rect 219 7608 231 7642
rect 1607 7608 1619 7642
rect 132 7594 178 7606
rect 219 7602 1619 7608
rect 132 7560 138 7594
rect 172 7560 178 7594
rect 132 7548 178 7560
rect 219 7546 1619 7552
rect 219 7512 231 7546
rect 1607 7512 1619 7546
rect 219 7506 1619 7512
rect 1660 7498 1706 7510
rect 1660 7464 1666 7498
rect 1700 7464 1706 7498
rect 219 7450 1619 7456
rect 1660 7452 1706 7464
rect 219 7416 231 7450
rect 1607 7416 1619 7450
rect 132 7402 178 7414
rect 219 7410 1619 7416
rect 132 7368 138 7402
rect 172 7368 178 7402
rect 132 7356 178 7368
rect 219 7354 1619 7360
rect 219 7320 231 7354
rect 1607 7320 1619 7354
rect 219 7314 1619 7320
rect 1660 7306 1706 7318
rect 1660 7272 1666 7306
rect 1700 7272 1706 7306
rect 219 7258 1619 7264
rect 1660 7260 1706 7272
rect 219 7224 231 7258
rect 1607 7224 1619 7258
rect 132 7210 178 7222
rect 219 7218 1619 7224
rect 132 7176 138 7210
rect 172 7176 178 7210
rect 132 7164 178 7176
rect 219 7162 1619 7168
rect 219 7128 231 7162
rect 1607 7128 1619 7162
rect 219 7122 1619 7128
rect 1660 7114 1706 7126
rect 1660 7080 1666 7114
rect 1700 7080 1706 7114
rect 219 7066 1619 7072
rect 1660 7068 1706 7080
rect 219 7032 231 7066
rect 1607 7032 1619 7066
rect 132 7018 178 7030
rect 219 7026 1619 7032
rect 132 6984 138 7018
rect 172 6984 178 7018
rect 132 6972 178 6984
rect 219 6970 1619 6976
rect 219 6936 231 6970
rect 1607 6936 1619 6970
rect 219 6930 1619 6936
rect 1660 6922 1706 6934
rect 1660 6888 1666 6922
rect 1700 6888 1706 6922
rect 219 6874 1619 6880
rect 1660 6876 1706 6888
rect 219 6840 231 6874
rect 1607 6840 1619 6874
rect 132 6826 178 6838
rect 219 6834 1619 6840
rect 132 6792 138 6826
rect 172 6792 178 6826
rect 132 6780 178 6792
rect 219 6778 1619 6784
rect 219 6744 231 6778
rect 1607 6744 1619 6778
rect 219 6738 1619 6744
rect 1660 6730 1706 6742
rect 1660 6696 1666 6730
rect 1700 6696 1706 6730
rect 219 6682 1619 6688
rect 1660 6684 1706 6696
rect 219 6648 231 6682
rect 1607 6648 1619 6682
rect 132 6634 178 6646
rect 219 6642 1619 6648
rect 132 6600 138 6634
rect 172 6600 178 6634
rect 132 6588 178 6600
rect 219 6586 1619 6592
rect 219 6552 231 6586
rect 1607 6552 1619 6586
rect 219 6546 1619 6552
rect 1660 6538 1706 6550
rect 1660 6504 1666 6538
rect 1700 6504 1706 6538
rect 219 6490 1619 6496
rect 1660 6492 1706 6504
rect 219 6456 231 6490
rect 1607 6456 1619 6490
rect 132 6442 178 6454
rect 219 6450 1619 6456
rect 132 6408 138 6442
rect 172 6408 178 6442
rect 132 6396 178 6408
rect 219 6394 1619 6400
rect 219 6360 231 6394
rect 1607 6360 1619 6394
rect 219 6354 1619 6360
rect 1660 6346 1706 6358
rect 1660 6312 1666 6346
rect 1700 6312 1706 6346
rect 219 6298 1619 6304
rect 1660 6300 1706 6312
rect 219 6264 231 6298
rect 1607 6264 1619 6298
rect 132 6250 178 6262
rect 219 6258 1619 6264
rect 132 6216 138 6250
rect 172 6216 178 6250
rect 132 6204 178 6216
rect 219 6202 1619 6208
rect 219 6168 231 6202
rect 1607 6168 1619 6202
rect 219 6162 1619 6168
rect 1660 6154 1706 6166
rect 1660 6120 1666 6154
rect 1700 6120 1706 6154
rect 219 6106 1619 6112
rect 1660 6108 1706 6120
rect 219 6072 231 6106
rect 1607 6072 1619 6106
rect 132 6058 178 6070
rect 219 6066 1619 6072
rect 132 6024 138 6058
rect 172 6024 178 6058
rect 132 6012 178 6024
rect 219 6010 1619 6016
rect 219 5976 231 6010
rect 1607 5976 1619 6010
rect 219 5970 1619 5976
rect 1660 5962 1706 5974
rect 1660 5928 1666 5962
rect 1700 5928 1706 5962
rect 219 5914 1619 5920
rect 1660 5916 1706 5928
rect 219 5880 231 5914
rect 1607 5880 1619 5914
rect 132 5866 178 5878
rect 219 5874 1619 5880
rect 132 5832 138 5866
rect 172 5832 178 5866
rect 132 5820 178 5832
rect 219 5818 1619 5824
rect 219 5784 231 5818
rect 1607 5784 1619 5818
rect 219 5778 1619 5784
rect 1660 5770 1706 5782
rect 1660 5736 1666 5770
rect 1700 5736 1706 5770
rect 219 5722 1619 5728
rect 1660 5724 1706 5736
rect 219 5688 231 5722
rect 1607 5688 1619 5722
rect 132 5674 178 5686
rect 219 5682 1619 5688
rect 132 5640 138 5674
rect 172 5640 178 5674
rect 132 5628 178 5640
rect 219 5626 1619 5632
rect 219 5592 231 5626
rect 1607 5592 1619 5626
rect 219 5586 1619 5592
rect 1660 5578 1706 5590
rect 1660 5544 1666 5578
rect 1700 5544 1706 5578
rect 219 5530 1619 5536
rect 1660 5532 1706 5544
rect 219 5496 231 5530
rect 1607 5496 1619 5530
rect 132 5482 178 5494
rect 219 5490 1619 5496
rect 132 5448 138 5482
rect 172 5448 178 5482
rect 132 5436 178 5448
rect 219 5434 1619 5440
rect 219 5400 231 5434
rect 1607 5400 1619 5434
rect 219 5394 1619 5400
rect 1660 5386 1706 5398
rect 1660 5352 1666 5386
rect 1700 5352 1706 5386
rect 219 5338 1619 5344
rect 1660 5340 1706 5352
rect 219 5304 231 5338
rect 1607 5304 1619 5338
rect 132 5290 178 5302
rect 219 5298 1619 5304
rect 132 5256 138 5290
rect 172 5256 178 5290
rect 132 5244 178 5256
rect 219 5242 1619 5248
rect 219 5208 231 5242
rect 1607 5208 1619 5242
rect 219 5202 1619 5208
rect 1660 5194 1706 5206
rect 1660 5160 1666 5194
rect 1700 5160 1706 5194
rect 219 5146 1619 5152
rect 1660 5148 1706 5160
rect 219 5112 231 5146
rect 1607 5112 1619 5146
rect 132 5098 178 5110
rect 219 5106 1619 5112
rect 132 5064 138 5098
rect 172 5064 178 5098
rect 132 5052 178 5064
rect 219 5050 1619 5056
rect 219 5016 231 5050
rect 1607 5016 1619 5050
rect 219 5010 1619 5016
rect 1660 5002 1706 5014
rect 1660 4968 1666 5002
rect 1700 4968 1706 5002
rect 219 4954 1619 4960
rect 1660 4956 1706 4968
rect 219 4920 231 4954
rect 1607 4920 1619 4954
rect 132 4906 178 4918
rect 219 4914 1619 4920
rect 132 4872 138 4906
rect 172 4872 178 4906
rect 132 4860 178 4872
rect 219 4858 1619 4864
rect 219 4824 231 4858
rect 1607 4824 1619 4858
rect 219 4818 1619 4824
rect 1660 4810 1706 4822
rect 1660 4776 1666 4810
rect 1700 4776 1706 4810
rect 219 4762 1619 4768
rect 1660 4764 1706 4776
rect 219 4728 231 4762
rect 1607 4728 1619 4762
rect 132 4714 178 4726
rect 219 4722 1619 4728
rect 132 4680 138 4714
rect 172 4680 178 4714
rect 132 4668 178 4680
rect 219 4666 1619 4672
rect 219 4632 231 4666
rect 1607 4632 1619 4666
rect 219 4626 1619 4632
rect 1660 4618 1706 4630
rect 1660 4584 1666 4618
rect 1700 4584 1706 4618
rect 219 4570 1619 4576
rect 1660 4572 1706 4584
rect 219 4536 231 4570
rect 1607 4536 1619 4570
rect 132 4522 178 4534
rect 219 4530 1619 4536
rect 132 4488 138 4522
rect 172 4488 178 4522
rect 132 4476 178 4488
rect 219 4474 1619 4480
rect 219 4440 231 4474
rect 1607 4440 1619 4474
rect 219 4434 1619 4440
rect 1660 4426 1706 4438
rect 1660 4392 1666 4426
rect 1700 4392 1706 4426
rect 219 4378 1619 4384
rect 1660 4380 1706 4392
rect 219 4344 231 4378
rect 1607 4344 1619 4378
rect 132 4330 178 4342
rect 219 4338 1619 4344
rect 132 4296 138 4330
rect 172 4296 178 4330
rect 132 4284 178 4296
rect 219 4282 1619 4288
rect 219 4248 231 4282
rect 1607 4248 1619 4282
rect 219 4242 1619 4248
rect 1660 4234 1706 4246
rect 1660 4200 1666 4234
rect 1700 4200 1706 4234
rect 219 4186 1619 4192
rect 1660 4188 1706 4200
rect 219 4152 231 4186
rect 1607 4152 1619 4186
rect 132 4138 178 4150
rect 219 4146 1619 4152
rect 132 4104 138 4138
rect 172 4104 178 4138
rect 132 4092 178 4104
rect 219 4090 1619 4096
rect 219 4056 231 4090
rect 1607 4056 1619 4090
rect 219 4050 1619 4056
rect 1660 4042 1706 4054
rect 1660 4008 1666 4042
rect 1700 4008 1706 4042
rect 219 3994 1619 4000
rect 1660 3996 1706 4008
rect 219 3960 231 3994
rect 1607 3960 1619 3994
rect 132 3946 178 3958
rect 219 3954 1619 3960
rect 132 3912 138 3946
rect 172 3912 178 3946
rect 132 3900 178 3912
rect 219 3898 1619 3904
rect 219 3864 231 3898
rect 1607 3864 1619 3898
rect 219 3858 1619 3864
rect 1660 3850 1706 3862
rect 1660 3816 1666 3850
rect 1700 3816 1706 3850
rect 219 3802 1619 3808
rect 1660 3804 1706 3816
rect 219 3768 231 3802
rect 1607 3768 1619 3802
rect 132 3754 178 3766
rect 219 3762 1619 3768
rect 132 3720 138 3754
rect 172 3720 178 3754
rect 132 3708 178 3720
rect 219 3706 1619 3712
rect 219 3672 231 3706
rect 1607 3672 1619 3706
rect 219 3666 1619 3672
rect 1660 3658 1706 3670
rect 1660 3624 1666 3658
rect 1700 3624 1706 3658
rect 219 3610 1619 3616
rect 1660 3612 1706 3624
rect 219 3576 231 3610
rect 1607 3576 1619 3610
rect 132 3562 178 3574
rect 219 3570 1619 3576
rect 132 3528 138 3562
rect 172 3528 178 3562
rect 132 3516 178 3528
rect 219 3514 1619 3520
rect 219 3480 231 3514
rect 1607 3480 1619 3514
rect 219 3474 1619 3480
rect 1660 3466 1706 3478
rect 1660 3432 1666 3466
rect 1700 3432 1706 3466
rect 219 3418 1619 3424
rect 1660 3420 1706 3432
rect 219 3384 231 3418
rect 1607 3384 1619 3418
rect 132 3370 178 3382
rect 219 3378 1619 3384
rect 132 3336 138 3370
rect 172 3336 178 3370
rect 132 3324 178 3336
rect 219 3322 1619 3328
rect 219 3288 231 3322
rect 1607 3288 1619 3322
rect 219 3282 1619 3288
rect 1660 3274 1706 3286
rect 1660 3240 1666 3274
rect 1700 3240 1706 3274
rect 219 3226 1619 3232
rect 1660 3228 1706 3240
rect 219 3192 231 3226
rect 1607 3192 1619 3226
rect 132 3178 178 3190
rect 219 3186 1619 3192
rect 132 3144 138 3178
rect 172 3144 178 3178
rect 132 3132 178 3144
rect 219 3130 1619 3136
rect 219 3096 231 3130
rect 1607 3096 1619 3130
rect 219 3090 1619 3096
rect 1660 3082 1706 3094
rect 1660 3048 1666 3082
rect 1700 3048 1706 3082
rect 219 3034 1619 3040
rect 1660 3036 1706 3048
rect 219 3000 231 3034
rect 1607 3000 1619 3034
rect 132 2986 178 2998
rect 219 2994 1619 3000
rect 132 2952 138 2986
rect 172 2952 178 2986
rect 132 2940 178 2952
rect 219 2938 1619 2944
rect 219 2904 231 2938
rect 1607 2904 1619 2938
rect 219 2898 1619 2904
rect 1660 2890 1706 2902
rect 1660 2856 1666 2890
rect 1700 2856 1706 2890
rect 219 2842 1619 2848
rect 1660 2844 1706 2856
rect 219 2808 231 2842
rect 1607 2808 1619 2842
rect 132 2794 178 2806
rect 219 2802 1619 2808
rect 132 2760 138 2794
rect 172 2760 178 2794
rect 132 2748 178 2760
rect 219 2746 1619 2752
rect 219 2712 231 2746
rect 1607 2712 1619 2746
rect 219 2706 1619 2712
rect 1660 2698 1706 2710
rect 1660 2664 1666 2698
rect 1700 2664 1706 2698
rect 219 2650 1619 2656
rect 1660 2652 1706 2664
rect 219 2616 231 2650
rect 1607 2616 1619 2650
rect 132 2602 178 2614
rect 219 2610 1619 2616
rect 132 2568 138 2602
rect 172 2568 178 2602
rect 132 2556 178 2568
rect 219 2554 1619 2560
rect 219 2520 231 2554
rect 1607 2520 1619 2554
rect 219 2514 1619 2520
rect 1660 2506 1706 2518
rect 1660 2472 1666 2506
rect 1700 2472 1706 2506
rect 219 2458 1619 2464
rect 1660 2460 1706 2472
rect 219 2424 231 2458
rect 1607 2424 1619 2458
rect 132 2410 178 2422
rect 219 2418 1619 2424
rect 132 2376 138 2410
rect 172 2376 178 2410
rect 132 2364 178 2376
rect 219 2362 1619 2368
rect 219 2328 231 2362
rect 1607 2328 1619 2362
rect 219 2322 1619 2328
rect 1660 2314 1706 2326
rect 1660 2280 1666 2314
rect 1700 2280 1706 2314
rect 219 2266 1619 2272
rect 1660 2268 1706 2280
rect 219 2232 231 2266
rect 1607 2232 1619 2266
rect 132 2218 178 2230
rect 219 2226 1619 2232
rect 132 2184 138 2218
rect 172 2184 178 2218
rect 132 2172 178 2184
rect 219 2170 1619 2176
rect 219 2136 231 2170
rect 1607 2136 1619 2170
rect 219 2130 1619 2136
rect 1660 2122 1706 2134
rect 1660 2088 1666 2122
rect 1700 2088 1706 2122
rect 219 2074 1619 2080
rect 1660 2076 1706 2088
rect 219 2040 231 2074
rect 1607 2040 1619 2074
rect 132 2026 178 2038
rect 219 2034 1619 2040
rect 132 1992 138 2026
rect 172 1992 178 2026
rect 132 1980 178 1992
rect 219 1978 1619 1984
rect 219 1944 231 1978
rect 1607 1944 1619 1978
rect 219 1938 1619 1944
rect 1660 1930 1706 1942
rect 1660 1896 1666 1930
rect 1700 1896 1706 1930
rect 219 1882 1619 1888
rect 1660 1884 1706 1896
rect 219 1848 231 1882
rect 1607 1848 1619 1882
rect 132 1834 178 1846
rect 219 1842 1619 1848
rect 132 1800 138 1834
rect 172 1800 178 1834
rect 132 1788 178 1800
rect 219 1786 1619 1792
rect 219 1752 231 1786
rect 1607 1752 1619 1786
rect 219 1746 1619 1752
rect 1660 1738 1706 1750
rect 1660 1704 1666 1738
rect 1700 1704 1706 1738
rect 219 1690 1619 1696
rect 1660 1692 1706 1704
rect 219 1656 231 1690
rect 1607 1656 1619 1690
rect 132 1642 178 1654
rect 219 1650 1619 1656
rect 132 1608 138 1642
rect 172 1608 178 1642
rect 132 1596 178 1608
rect 219 1594 1619 1600
rect 219 1560 231 1594
rect 1607 1560 1619 1594
rect 219 1554 1619 1560
rect 1660 1546 1706 1558
rect 1660 1512 1666 1546
rect 1700 1512 1706 1546
rect 219 1498 1619 1504
rect 1660 1500 1706 1512
rect 219 1464 231 1498
rect 1607 1464 1619 1498
rect 132 1450 178 1462
rect 219 1458 1619 1464
rect 132 1416 138 1450
rect 172 1416 178 1450
rect 132 1404 178 1416
rect 219 1402 1619 1408
rect 219 1368 231 1402
rect 1607 1368 1619 1402
rect 219 1362 1619 1368
rect 1660 1354 1706 1366
rect 1660 1320 1666 1354
rect 1700 1320 1706 1354
rect 219 1306 1619 1312
rect 1660 1308 1706 1320
rect 219 1272 231 1306
rect 1607 1272 1619 1306
rect 132 1258 178 1270
rect 219 1266 1619 1272
rect 132 1224 138 1258
rect 172 1224 178 1258
rect 132 1212 178 1224
rect 219 1210 1619 1216
rect 219 1176 231 1210
rect 1607 1176 1619 1210
rect 219 1170 1619 1176
rect 1660 1162 1706 1174
rect 1660 1128 1666 1162
rect 1700 1128 1706 1162
rect 219 1114 1619 1120
rect 1660 1116 1706 1128
rect 219 1080 231 1114
rect 1607 1080 1619 1114
rect 132 1066 178 1078
rect 219 1074 1619 1080
rect 132 1032 138 1066
rect 172 1032 178 1066
rect 132 1020 178 1032
rect 219 1018 1619 1024
rect 219 984 231 1018
rect 1607 984 1619 1018
rect 219 978 1619 984
rect 1660 970 1706 982
rect 1660 936 1666 970
rect 1700 936 1706 970
rect 219 922 1619 928
rect 1660 924 1706 936
rect 219 888 231 922
rect 1607 888 1619 922
rect 132 874 178 886
rect 219 882 1619 888
rect 132 840 138 874
rect 172 840 178 874
rect 132 828 178 840
rect 219 826 1619 832
rect 219 792 231 826
rect 1607 792 1619 826
rect 219 786 1619 792
rect 1660 778 1706 790
rect 1660 744 1666 778
rect 1700 744 1706 778
rect 219 730 1619 736
rect 1660 732 1706 744
rect 219 696 231 730
rect 1607 696 1619 730
rect 219 690 1619 696
<< metal4 >>
rect 0 22204 1840 22304
rect 0 0 240 22000
rect 340 0 870 22000
rect 970 0 1500 22000
rect 1600 0 1840 22000
<< labels >>
rlabel metal4 0 0 240 22000 1 VGND
port 1 n ground input
rlabel metal4 1600 0 1840 22000 1 VGND
port 1 n ground input
rlabel metal4 340 0 870 22000 1 VPWR
port 2 n power input
rlabel metal4 970 0 1500 22000 1 GPWR
port 3 n power output
rlabel metal4 0 22204 1840 22304 1 ctrl
port 4 n signal input
<< end >>
