magic
tech sky130A
magscale 1 2
timestamp 1697722671
<< metal1 >>
rect -10593 -60 -10527 -50
rect -10593 -576 -10527 -566
rect -10401 -60 -10335 -50
rect -10401 -576 -10335 -566
rect -10209 -60 -10143 -50
rect -10209 -576 -10143 -566
rect -10017 -60 -9951 -50
rect -10017 -576 -9951 -566
rect -9825 -60 -9759 -50
rect -9825 -576 -9759 -566
rect -9633 -60 -9567 -50
rect -9633 -576 -9567 -566
rect -9441 -60 -9375 -50
rect -9441 -576 -9375 -566
rect -9249 -60 -9183 -50
rect -9249 -576 -9183 -566
rect -9057 -60 -8991 -50
rect -9057 -576 -8991 -566
rect -8865 -60 -8799 -50
rect -8865 -576 -8799 -566
rect -8673 -60 -8607 -50
rect -8673 -576 -8607 -566
rect -8481 -60 -8415 -50
rect -8481 -576 -8415 -566
rect -8289 -60 -8223 -50
rect -8289 -576 -8223 -566
rect -8097 -60 -8031 -50
rect -8097 -576 -8031 -566
rect -7905 -60 -7839 -50
rect -7905 -576 -7839 -566
rect -7713 -60 -7647 -50
rect -7713 -576 -7647 -566
rect -7521 -60 -7455 -50
rect -7521 -576 -7455 -566
rect -7329 -60 -7263 -50
rect -7329 -576 -7263 -566
rect -7137 -60 -7071 -50
rect -7137 -576 -7071 -566
rect -6945 -60 -6879 -50
rect -6945 -576 -6879 -566
rect -6753 -60 -6687 -50
rect -6753 -576 -6687 -566
rect -6561 -60 -6495 -50
rect -6561 -576 -6495 -566
rect -6369 -60 -6303 -50
rect -6369 -576 -6303 -566
rect -6177 -60 -6111 -50
rect -6177 -576 -6111 -566
rect -5985 -60 -5919 -50
rect -5985 -576 -5919 -566
rect -5793 -60 -5727 -50
rect -5793 -576 -5727 -566
rect -5601 -60 -5535 -50
rect -5601 -576 -5535 -566
rect -5409 -60 -5343 -50
rect -5409 -576 -5343 -566
rect -5217 -60 -5151 -50
rect -5217 -576 -5151 -566
rect -5025 -60 -4959 -50
rect -5025 -576 -4959 -566
rect -4833 -60 -4767 -50
rect -4833 -576 -4767 -566
rect -4641 -60 -4575 -50
rect -4641 -576 -4575 -566
rect -4449 -60 -4383 -50
rect -4449 -576 -4383 -566
rect -4257 -60 -4191 -50
rect -4257 -576 -4191 -566
rect -4065 -60 -3999 -50
rect -4065 -576 -3999 -566
rect -3873 -60 -3807 -50
rect -3873 -576 -3807 -566
rect -3681 -60 -3615 -50
rect -3681 -576 -3615 -566
rect -3489 -60 -3423 -50
rect -3489 -576 -3423 -566
rect -3297 -60 -3231 -50
rect -3297 -576 -3231 -566
rect -3105 -60 -3039 -50
rect -3105 -576 -3039 -566
rect -2913 -60 -2847 -50
rect -2913 -576 -2847 -566
rect -2721 -60 -2655 -50
rect -2721 -576 -2655 -566
rect -2529 -60 -2463 -50
rect -2529 -576 -2463 -566
rect -2337 -60 -2271 -50
rect -2337 -576 -2271 -566
rect -2145 -60 -2079 -50
rect -2145 -576 -2079 -566
rect -1953 -60 -1887 -50
rect -1953 -576 -1887 -566
rect -1761 -60 -1695 -50
rect -1761 -576 -1695 -566
rect -1569 -60 -1503 -50
rect -1569 -576 -1503 -566
rect -1377 -60 -1311 -50
rect -1377 -576 -1311 -566
rect -1185 -60 -1119 -50
rect -1185 -576 -1119 -566
rect -993 -60 -927 -50
rect -993 -576 -927 -566
rect -801 -60 -735 -50
rect -801 -576 -735 -566
rect -609 -60 -543 -50
rect -609 -576 -543 -566
rect -417 -60 -351 -50
rect -417 -576 -351 -566
rect -225 -60 -159 -50
rect -225 -576 -159 -566
rect -33 -60 33 -50
rect -33 -576 33 -566
rect 159 -60 225 -50
rect 159 -576 225 -566
rect 351 -60 417 -50
rect 351 -576 417 -566
rect 543 -60 609 -50
rect 543 -576 609 -566
rect 735 -60 801 -50
rect 735 -576 801 -566
rect 927 -60 993 -50
rect 927 -576 993 -566
rect 1119 -60 1185 -50
rect 1119 -576 1185 -566
rect 1311 -60 1377 -50
rect 1311 -576 1377 -566
rect 1503 -60 1569 -50
rect 1503 -576 1569 -566
rect 1695 -60 1761 -50
rect 1695 -576 1761 -566
rect 1887 -60 1953 -50
rect 1887 -576 1953 -566
rect 2079 -60 2145 -50
rect 2079 -576 2145 -566
rect 2271 -60 2337 -50
rect 2271 -576 2337 -566
rect 2463 -60 2529 -50
rect 2463 -576 2529 -566
rect 2655 -60 2721 -50
rect 2655 -576 2721 -566
rect 2847 -60 2913 -50
rect 2847 -576 2913 -566
rect 3039 -60 3105 -50
rect 3039 -576 3105 -566
rect 3231 -60 3297 -50
rect 3231 -576 3297 -566
rect 3423 -60 3489 -50
rect 3423 -576 3489 -566
rect 3615 -60 3681 -50
rect 3615 -576 3681 -566
rect 3807 -60 3873 -50
rect 3807 -576 3873 -566
rect 3999 -60 4065 -50
rect 3999 -576 4065 -566
rect 4191 -60 4257 -50
rect 4191 -576 4257 -566
rect 4383 -60 4449 -50
rect 4383 -576 4449 -566
rect 4575 -60 4641 -50
rect 4575 -576 4641 -566
rect 4767 -60 4833 -50
rect 4767 -576 4833 -566
rect 4959 -60 5025 -50
rect 4959 -576 5025 -566
rect 5151 -60 5217 -50
rect 5151 -576 5217 -566
rect 5343 -60 5409 -50
rect 5343 -576 5409 -566
rect 5535 -60 5601 -50
rect 5535 -576 5601 -566
rect 5727 -60 5793 -50
rect 5727 -576 5793 -566
rect 5919 -60 5985 -50
rect 5919 -576 5985 -566
rect 6111 -60 6177 -50
rect 6111 -576 6177 -566
rect 6303 -60 6369 -50
rect 6303 -576 6369 -566
rect 6495 -60 6561 -50
rect 6495 -576 6561 -566
rect 6687 -60 6753 -50
rect 6687 -576 6753 -566
rect 6879 -60 6945 -50
rect 6879 -576 6945 -566
rect 7071 -60 7137 -50
rect 7071 -576 7137 -566
rect 7263 -60 7329 -50
rect 7263 -576 7329 -566
rect 7455 -60 7521 -50
rect 7455 -576 7521 -566
rect 7647 -60 7713 -50
rect 7647 -576 7713 -566
rect 7839 -60 7905 -50
rect 7839 -576 7905 -566
rect 8031 -60 8097 -50
rect 8031 -576 8097 -566
rect 8223 -60 8289 -50
rect 8223 -576 8289 -566
rect 8415 -60 8481 -50
rect 8415 -576 8481 -566
rect 8607 -60 8673 -50
rect 8607 -576 8673 -566
rect 8799 -60 8865 -50
rect 8799 -576 8865 -566
rect 8991 -60 9057 -50
rect 8991 -576 9057 -566
rect 9183 -60 9249 -50
rect 9183 -576 9249 -566
rect 9375 -60 9441 -50
rect 9375 -576 9441 -566
rect 9567 -60 9633 -50
rect 9567 -576 9633 -566
rect 9759 -60 9825 -50
rect 9759 -576 9825 -566
rect 9951 -60 10017 -50
rect 9951 -576 10017 -566
rect 10143 -60 10209 -50
rect 10143 -576 10209 -566
rect 10335 -60 10401 -50
rect 10335 -576 10401 -566
rect 10527 -60 10593 -50
rect 10527 -576 10593 -566
<< via1 >>
rect -10593 -566 -10527 -60
rect -10401 -566 -10335 -60
rect -10209 -566 -10143 -60
rect -10017 -566 -9951 -60
rect -9825 -566 -9759 -60
rect -9633 -566 -9567 -60
rect -9441 -566 -9375 -60
rect -9249 -566 -9183 -60
rect -9057 -566 -8991 -60
rect -8865 -566 -8799 -60
rect -8673 -566 -8607 -60
rect -8481 -566 -8415 -60
rect -8289 -566 -8223 -60
rect -8097 -566 -8031 -60
rect -7905 -566 -7839 -60
rect -7713 -566 -7647 -60
rect -7521 -566 -7455 -60
rect -7329 -566 -7263 -60
rect -7137 -566 -7071 -60
rect -6945 -566 -6879 -60
rect -6753 -566 -6687 -60
rect -6561 -566 -6495 -60
rect -6369 -566 -6303 -60
rect -6177 -566 -6111 -60
rect -5985 -566 -5919 -60
rect -5793 -566 -5727 -60
rect -5601 -566 -5535 -60
rect -5409 -566 -5343 -60
rect -5217 -566 -5151 -60
rect -5025 -566 -4959 -60
rect -4833 -566 -4767 -60
rect -4641 -566 -4575 -60
rect -4449 -566 -4383 -60
rect -4257 -566 -4191 -60
rect -4065 -566 -3999 -60
rect -3873 -566 -3807 -60
rect -3681 -566 -3615 -60
rect -3489 -566 -3423 -60
rect -3297 -566 -3231 -60
rect -3105 -566 -3039 -60
rect -2913 -566 -2847 -60
rect -2721 -566 -2655 -60
rect -2529 -566 -2463 -60
rect -2337 -566 -2271 -60
rect -2145 -566 -2079 -60
rect -1953 -566 -1887 -60
rect -1761 -566 -1695 -60
rect -1569 -566 -1503 -60
rect -1377 -566 -1311 -60
rect -1185 -566 -1119 -60
rect -993 -566 -927 -60
rect -801 -566 -735 -60
rect -609 -566 -543 -60
rect -417 -566 -351 -60
rect -225 -566 -159 -60
rect -33 -566 33 -60
rect 159 -566 225 -60
rect 351 -566 417 -60
rect 543 -566 609 -60
rect 735 -566 801 -60
rect 927 -566 993 -60
rect 1119 -566 1185 -60
rect 1311 -566 1377 -60
rect 1503 -566 1569 -60
rect 1695 -566 1761 -60
rect 1887 -566 1953 -60
rect 2079 -566 2145 -60
rect 2271 -566 2337 -60
rect 2463 -566 2529 -60
rect 2655 -566 2721 -60
rect 2847 -566 2913 -60
rect 3039 -566 3105 -60
rect 3231 -566 3297 -60
rect 3423 -566 3489 -60
rect 3615 -566 3681 -60
rect 3807 -566 3873 -60
rect 3999 -566 4065 -60
rect 4191 -566 4257 -60
rect 4383 -566 4449 -60
rect 4575 -566 4641 -60
rect 4767 -566 4833 -60
rect 4959 -566 5025 -60
rect 5151 -566 5217 -60
rect 5343 -566 5409 -60
rect 5535 -566 5601 -60
rect 5727 -566 5793 -60
rect 5919 -566 5985 -60
rect 6111 -566 6177 -60
rect 6303 -566 6369 -60
rect 6495 -566 6561 -60
rect 6687 -566 6753 -60
rect 6879 -566 6945 -60
rect 7071 -566 7137 -60
rect 7263 -566 7329 -60
rect 7455 -566 7521 -60
rect 7647 -566 7713 -60
rect 7839 -566 7905 -60
rect 8031 -566 8097 -60
rect 8223 -566 8289 -60
rect 8415 -566 8481 -60
rect 8607 -566 8673 -60
rect 8799 -566 8865 -60
rect 8991 -566 9057 -60
rect 9183 -566 9249 -60
rect 9375 -566 9441 -60
rect 9567 -566 9633 -60
rect 9759 -566 9825 -60
rect 9951 -566 10017 -60
rect 10143 -566 10209 -60
rect 10335 -566 10401 -60
rect 10527 -566 10593 -60
<< metal2 >>
rect -10603 -60 -10517 -50
rect -10603 -566 -10593 -60
rect -10527 -566 -10517 -60
rect -10603 -576 -10517 -566
rect -10411 -60 -10325 -50
rect -10411 -566 -10401 -60
rect -10335 -566 -10325 -60
rect -10411 -576 -10325 -566
rect -10219 -60 -10133 -50
rect -10219 -566 -10209 -60
rect -10143 -566 -10133 -60
rect -10219 -576 -10133 -566
rect -10027 -60 -9941 -50
rect -10027 -566 -10017 -60
rect -9951 -566 -9941 -60
rect -10027 -576 -9941 -566
rect -9835 -60 -9749 -50
rect -9835 -566 -9825 -60
rect -9759 -566 -9749 -60
rect -9835 -576 -9749 -566
rect -9643 -60 -9557 -50
rect -9643 -566 -9633 -60
rect -9567 -566 -9557 -60
rect -9643 -576 -9557 -566
rect -9451 -60 -9365 -50
rect -9451 -566 -9441 -60
rect -9375 -566 -9365 -60
rect -9451 -576 -9365 -566
rect -9259 -60 -9173 -50
rect -9259 -566 -9249 -60
rect -9183 -566 -9173 -60
rect -9259 -576 -9173 -566
rect -9067 -60 -8981 -50
rect -9067 -566 -9057 -60
rect -8991 -566 -8981 -60
rect -9067 -576 -8981 -566
rect -8875 -60 -8789 -50
rect -8875 -566 -8865 -60
rect -8799 -566 -8789 -60
rect -8875 -576 -8789 -566
rect -8683 -60 -8597 -50
rect -8683 -566 -8673 -60
rect -8607 -566 -8597 -60
rect -8683 -576 -8597 -566
rect -8491 -60 -8405 -50
rect -8491 -566 -8481 -60
rect -8415 -566 -8405 -60
rect -8491 -576 -8405 -566
rect -8299 -60 -8213 -50
rect -8299 -566 -8289 -60
rect -8223 -566 -8213 -60
rect -8299 -576 -8213 -566
rect -8107 -60 -8021 -50
rect -8107 -566 -8097 -60
rect -8031 -566 -8021 -60
rect -8107 -576 -8021 -566
rect -7915 -60 -7829 -50
rect -7915 -566 -7905 -60
rect -7839 -566 -7829 -60
rect -7915 -576 -7829 -566
rect -7723 -60 -7637 -50
rect -7723 -566 -7713 -60
rect -7647 -566 -7637 -60
rect -7723 -576 -7637 -566
rect -7531 -60 -7445 -50
rect -7531 -566 -7521 -60
rect -7455 -566 -7445 -60
rect -7531 -576 -7445 -566
rect -7339 -60 -7253 -50
rect -7339 -566 -7329 -60
rect -7263 -566 -7253 -60
rect -7339 -576 -7253 -566
rect -7147 -60 -7061 -50
rect -7147 -566 -7137 -60
rect -7071 -566 -7061 -60
rect -7147 -576 -7061 -566
rect -6955 -60 -6869 -50
rect -6955 -566 -6945 -60
rect -6879 -566 -6869 -60
rect -6955 -576 -6869 -566
rect -6763 -60 -6677 -50
rect -6763 -566 -6753 -60
rect -6687 -566 -6677 -60
rect -6763 -576 -6677 -566
rect -6571 -60 -6485 -50
rect -6571 -566 -6561 -60
rect -6495 -566 -6485 -60
rect -6571 -576 -6485 -566
rect -6379 -60 -6293 -50
rect -6379 -566 -6369 -60
rect -6303 -566 -6293 -60
rect -6379 -576 -6293 -566
rect -6187 -60 -6101 -50
rect -6187 -566 -6177 -60
rect -6111 -566 -6101 -60
rect -6187 -576 -6101 -566
rect -5995 -60 -5909 -50
rect -5995 -566 -5985 -60
rect -5919 -566 -5909 -60
rect -5995 -576 -5909 -566
rect -5803 -60 -5717 -50
rect -5803 -566 -5793 -60
rect -5727 -566 -5717 -60
rect -5803 -576 -5717 -566
rect -5611 -60 -5525 -50
rect -5611 -566 -5601 -60
rect -5535 -566 -5525 -60
rect -5611 -576 -5525 -566
rect -5419 -60 -5333 -50
rect -5419 -566 -5409 -60
rect -5343 -566 -5333 -60
rect -5419 -576 -5333 -566
rect -5227 -60 -5141 -50
rect -5227 -566 -5217 -60
rect -5151 -566 -5141 -60
rect -5227 -576 -5141 -566
rect -5035 -60 -4949 -50
rect -5035 -566 -5025 -60
rect -4959 -566 -4949 -60
rect -5035 -576 -4949 -566
rect -4843 -60 -4757 -50
rect -4843 -566 -4833 -60
rect -4767 -566 -4757 -60
rect -4843 -576 -4757 -566
rect -4651 -60 -4565 -50
rect -4651 -566 -4641 -60
rect -4575 -566 -4565 -60
rect -4651 -576 -4565 -566
rect -4459 -60 -4373 -50
rect -4459 -566 -4449 -60
rect -4383 -566 -4373 -60
rect -4459 -576 -4373 -566
rect -4267 -60 -4181 -50
rect -4267 -566 -4257 -60
rect -4191 -566 -4181 -60
rect -4267 -576 -4181 -566
rect -4075 -60 -3989 -50
rect -4075 -566 -4065 -60
rect -3999 -566 -3989 -60
rect -4075 -576 -3989 -566
rect -3883 -60 -3797 -50
rect -3883 -566 -3873 -60
rect -3807 -566 -3797 -60
rect -3883 -576 -3797 -566
rect -3691 -60 -3605 -50
rect -3691 -566 -3681 -60
rect -3615 -566 -3605 -60
rect -3691 -576 -3605 -566
rect -3499 -60 -3413 -50
rect -3499 -566 -3489 -60
rect -3423 -566 -3413 -60
rect -3499 -576 -3413 -566
rect -3307 -60 -3221 -50
rect -3307 -566 -3297 -60
rect -3231 -566 -3221 -60
rect -3307 -576 -3221 -566
rect -3115 -60 -3029 -50
rect -3115 -566 -3105 -60
rect -3039 -566 -3029 -60
rect -3115 -576 -3029 -566
rect -2923 -60 -2837 -50
rect -2923 -566 -2913 -60
rect -2847 -566 -2837 -60
rect -2923 -576 -2837 -566
rect -2731 -60 -2645 -50
rect -2731 -566 -2721 -60
rect -2655 -566 -2645 -60
rect -2731 -576 -2645 -566
rect -2539 -60 -2453 -50
rect -2539 -566 -2529 -60
rect -2463 -566 -2453 -60
rect -2539 -576 -2453 -566
rect -2347 -60 -2261 -50
rect -2347 -566 -2337 -60
rect -2271 -566 -2261 -60
rect -2347 -576 -2261 -566
rect -2155 -60 -2069 -50
rect -2155 -566 -2145 -60
rect -2079 -566 -2069 -60
rect -2155 -576 -2069 -566
rect -1963 -60 -1877 -50
rect -1963 -566 -1953 -60
rect -1887 -566 -1877 -60
rect -1963 -576 -1877 -566
rect -1771 -60 -1685 -50
rect -1771 -566 -1761 -60
rect -1695 -566 -1685 -60
rect -1771 -576 -1685 -566
rect -1579 -60 -1493 -50
rect -1579 -566 -1569 -60
rect -1503 -566 -1493 -60
rect -1579 -576 -1493 -566
rect -1387 -60 -1301 -50
rect -1387 -566 -1377 -60
rect -1311 -566 -1301 -60
rect -1387 -576 -1301 -566
rect -1195 -60 -1109 -50
rect -1195 -566 -1185 -60
rect -1119 -566 -1109 -60
rect -1195 -576 -1109 -566
rect -1003 -60 -917 -50
rect -1003 -566 -993 -60
rect -927 -566 -917 -60
rect -1003 -576 -917 -566
rect -811 -60 -725 -50
rect -811 -566 -801 -60
rect -735 -566 -725 -60
rect -811 -576 -725 -566
rect -619 -60 -533 -50
rect -619 -566 -609 -60
rect -543 -566 -533 -60
rect -619 -576 -533 -566
rect -427 -60 -341 -50
rect -427 -566 -417 -60
rect -351 -566 -341 -60
rect -427 -576 -341 -566
rect -235 -60 -149 -50
rect -235 -566 -225 -60
rect -159 -566 -149 -60
rect -235 -576 -149 -566
rect -43 -60 43 -50
rect -43 -566 -33 -60
rect 33 -566 43 -60
rect -43 -576 43 -566
rect 149 -60 235 -50
rect 149 -566 159 -60
rect 225 -566 235 -60
rect 149 -576 235 -566
rect 341 -60 427 -50
rect 341 -566 351 -60
rect 417 -566 427 -60
rect 341 -576 427 -566
rect 533 -60 619 -50
rect 533 -566 543 -60
rect 609 -566 619 -60
rect 533 -576 619 -566
rect 725 -60 811 -50
rect 725 -566 735 -60
rect 801 -566 811 -60
rect 725 -576 811 -566
rect 917 -60 1003 -50
rect 917 -566 927 -60
rect 993 -566 1003 -60
rect 917 -576 1003 -566
rect 1109 -60 1195 -50
rect 1109 -566 1119 -60
rect 1185 -566 1195 -60
rect 1109 -576 1195 -566
rect 1301 -60 1387 -50
rect 1301 -566 1311 -60
rect 1377 -566 1387 -60
rect 1301 -576 1387 -566
rect 1493 -60 1579 -50
rect 1493 -566 1503 -60
rect 1569 -566 1579 -60
rect 1493 -576 1579 -566
rect 1685 -60 1771 -50
rect 1685 -566 1695 -60
rect 1761 -566 1771 -60
rect 1685 -576 1771 -566
rect 1877 -60 1963 -50
rect 1877 -566 1887 -60
rect 1953 -566 1963 -60
rect 1877 -576 1963 -566
rect 2069 -60 2155 -50
rect 2069 -566 2079 -60
rect 2145 -566 2155 -60
rect 2069 -576 2155 -566
rect 2261 -60 2347 -50
rect 2261 -566 2271 -60
rect 2337 -566 2347 -60
rect 2261 -576 2347 -566
rect 2453 -60 2539 -50
rect 2453 -566 2463 -60
rect 2529 -566 2539 -60
rect 2453 -576 2539 -566
rect 2645 -60 2731 -50
rect 2645 -566 2655 -60
rect 2721 -566 2731 -60
rect 2645 -576 2731 -566
rect 2837 -60 2923 -50
rect 2837 -566 2847 -60
rect 2913 -566 2923 -60
rect 2837 -576 2923 -566
rect 3029 -60 3115 -50
rect 3029 -566 3039 -60
rect 3105 -566 3115 -60
rect 3029 -576 3115 -566
rect 3221 -60 3307 -50
rect 3221 -566 3231 -60
rect 3297 -566 3307 -60
rect 3221 -576 3307 -566
rect 3413 -60 3499 -50
rect 3413 -566 3423 -60
rect 3489 -566 3499 -60
rect 3413 -576 3499 -566
rect 3605 -60 3691 -50
rect 3605 -566 3615 -60
rect 3681 -566 3691 -60
rect 3605 -576 3691 -566
rect 3797 -60 3883 -50
rect 3797 -566 3807 -60
rect 3873 -566 3883 -60
rect 3797 -576 3883 -566
rect 3989 -60 4075 -50
rect 3989 -566 3999 -60
rect 4065 -566 4075 -60
rect 3989 -576 4075 -566
rect 4181 -60 4267 -50
rect 4181 -566 4191 -60
rect 4257 -566 4267 -60
rect 4181 -576 4267 -566
rect 4373 -60 4459 -50
rect 4373 -566 4383 -60
rect 4449 -566 4459 -60
rect 4373 -576 4459 -566
rect 4565 -60 4651 -50
rect 4565 -566 4575 -60
rect 4641 -566 4651 -60
rect 4565 -576 4651 -566
rect 4757 -60 4843 -50
rect 4757 -566 4767 -60
rect 4833 -566 4843 -60
rect 4757 -576 4843 -566
rect 4949 -60 5035 -50
rect 4949 -566 4959 -60
rect 5025 -566 5035 -60
rect 4949 -576 5035 -566
rect 5141 -60 5227 -50
rect 5141 -566 5151 -60
rect 5217 -566 5227 -60
rect 5141 -576 5227 -566
rect 5333 -60 5419 -50
rect 5333 -566 5343 -60
rect 5409 -566 5419 -60
rect 5333 -576 5419 -566
rect 5525 -60 5611 -50
rect 5525 -566 5535 -60
rect 5601 -566 5611 -60
rect 5525 -576 5611 -566
rect 5717 -60 5803 -50
rect 5717 -566 5727 -60
rect 5793 -566 5803 -60
rect 5717 -576 5803 -566
rect 5909 -60 5995 -50
rect 5909 -566 5919 -60
rect 5985 -566 5995 -60
rect 5909 -576 5995 -566
rect 6101 -60 6187 -50
rect 6101 -566 6111 -60
rect 6177 -566 6187 -60
rect 6101 -576 6187 -566
rect 6293 -60 6379 -50
rect 6293 -566 6303 -60
rect 6369 -566 6379 -60
rect 6293 -576 6379 -566
rect 6485 -60 6571 -50
rect 6485 -566 6495 -60
rect 6561 -566 6571 -60
rect 6485 -576 6571 -566
rect 6677 -60 6763 -50
rect 6677 -566 6687 -60
rect 6753 -566 6763 -60
rect 6677 -576 6763 -566
rect 6869 -60 6955 -50
rect 6869 -566 6879 -60
rect 6945 -566 6955 -60
rect 6869 -576 6955 -566
rect 7061 -60 7147 -50
rect 7061 -566 7071 -60
rect 7137 -566 7147 -60
rect 7061 -576 7147 -566
rect 7253 -60 7339 -50
rect 7253 -566 7263 -60
rect 7329 -566 7339 -60
rect 7253 -576 7339 -566
rect 7445 -60 7531 -50
rect 7445 -566 7455 -60
rect 7521 -566 7531 -60
rect 7445 -576 7531 -566
rect 7637 -60 7723 -50
rect 7637 -566 7647 -60
rect 7713 -566 7723 -60
rect 7637 -576 7723 -566
rect 7829 -60 7915 -50
rect 7829 -566 7839 -60
rect 7905 -566 7915 -60
rect 7829 -576 7915 -566
rect 8021 -60 8107 -50
rect 8021 -566 8031 -60
rect 8097 -566 8107 -60
rect 8021 -576 8107 -566
rect 8213 -60 8299 -50
rect 8213 -566 8223 -60
rect 8289 -566 8299 -60
rect 8213 -576 8299 -566
rect 8405 -60 8491 -50
rect 8405 -566 8415 -60
rect 8481 -566 8491 -60
rect 8405 -576 8491 -566
rect 8597 -60 8683 -50
rect 8597 -566 8607 -60
rect 8673 -566 8683 -60
rect 8597 -576 8683 -566
rect 8789 -60 8875 -50
rect 8789 -566 8799 -60
rect 8865 -566 8875 -60
rect 8789 -576 8875 -566
rect 8981 -60 9067 -50
rect 8981 -566 8991 -60
rect 9057 -566 9067 -60
rect 8981 -576 9067 -566
rect 9173 -60 9259 -50
rect 9173 -566 9183 -60
rect 9249 -566 9259 -60
rect 9173 -576 9259 -566
rect 9365 -60 9451 -50
rect 9365 -566 9375 -60
rect 9441 -566 9451 -60
rect 9365 -576 9451 -566
rect 9557 -60 9643 -50
rect 9557 -566 9567 -60
rect 9633 -566 9643 -60
rect 9557 -576 9643 -566
rect 9749 -60 9835 -50
rect 9749 -566 9759 -60
rect 9825 -566 9835 -60
rect 9749 -576 9835 -566
rect 9941 -60 10027 -50
rect 9941 -566 9951 -60
rect 10017 -566 10027 -60
rect 9941 -576 10027 -566
rect 10133 -60 10219 -50
rect 10133 -566 10143 -60
rect 10209 -566 10219 -60
rect 10133 -576 10219 -566
rect 10325 -60 10411 -50
rect 10325 -566 10335 -60
rect 10401 -566 10411 -60
rect 10325 -576 10411 -566
rect 10517 -60 10603 -50
rect 10517 -566 10527 -60
rect 10593 -566 10603 -60
rect 10517 -576 10603 -566
<< via2 >>
rect -10593 -566 -10527 -60
rect -10401 -566 -10335 -60
rect -10209 -566 -10143 -60
rect -10017 -566 -9951 -60
rect -9825 -566 -9759 -60
rect -9633 -566 -9567 -60
rect -9441 -566 -9375 -60
rect -9249 -566 -9183 -60
rect -9057 -566 -8991 -60
rect -8865 -566 -8799 -60
rect -8673 -566 -8607 -60
rect -8481 -566 -8415 -60
rect -8289 -566 -8223 -60
rect -8097 -566 -8031 -60
rect -7905 -566 -7839 -60
rect -7713 -566 -7647 -60
rect -7521 -566 -7455 -60
rect -7329 -566 -7263 -60
rect -7137 -566 -7071 -60
rect -6945 -566 -6879 -60
rect -6753 -566 -6687 -60
rect -6561 -566 -6495 -60
rect -6369 -566 -6303 -60
rect -6177 -566 -6111 -60
rect -5985 -566 -5919 -60
rect -5793 -566 -5727 -60
rect -5601 -566 -5535 -60
rect -5409 -566 -5343 -60
rect -5217 -566 -5151 -60
rect -5025 -566 -4959 -60
rect -4833 -566 -4767 -60
rect -4641 -566 -4575 -60
rect -4449 -566 -4383 -60
rect -4257 -566 -4191 -60
rect -4065 -566 -3999 -60
rect -3873 -566 -3807 -60
rect -3681 -566 -3615 -60
rect -3489 -566 -3423 -60
rect -3297 -566 -3231 -60
rect -3105 -566 -3039 -60
rect -2913 -566 -2847 -60
rect -2721 -566 -2655 -60
rect -2529 -566 -2463 -60
rect -2337 -566 -2271 -60
rect -2145 -566 -2079 -60
rect -1953 -566 -1887 -60
rect -1761 -566 -1695 -60
rect -1569 -566 -1503 -60
rect -1377 -566 -1311 -60
rect -1185 -566 -1119 -60
rect -993 -566 -927 -60
rect -801 -566 -735 -60
rect -609 -566 -543 -60
rect -417 -566 -351 -60
rect -225 -566 -159 -60
rect -33 -566 33 -60
rect 159 -566 225 -60
rect 351 -566 417 -60
rect 543 -566 609 -60
rect 735 -566 801 -60
rect 927 -566 993 -60
rect 1119 -566 1185 -60
rect 1311 -566 1377 -60
rect 1503 -566 1569 -60
rect 1695 -566 1761 -60
rect 1887 -566 1953 -60
rect 2079 -566 2145 -60
rect 2271 -566 2337 -60
rect 2463 -566 2529 -60
rect 2655 -566 2721 -60
rect 2847 -566 2913 -60
rect 3039 -566 3105 -60
rect 3231 -566 3297 -60
rect 3423 -566 3489 -60
rect 3615 -566 3681 -60
rect 3807 -566 3873 -60
rect 3999 -566 4065 -60
rect 4191 -566 4257 -60
rect 4383 -566 4449 -60
rect 4575 -566 4641 -60
rect 4767 -566 4833 -60
rect 4959 -566 5025 -60
rect 5151 -566 5217 -60
rect 5343 -566 5409 -60
rect 5535 -566 5601 -60
rect 5727 -566 5793 -60
rect 5919 -566 5985 -60
rect 6111 -566 6177 -60
rect 6303 -566 6369 -60
rect 6495 -566 6561 -60
rect 6687 -566 6753 -60
rect 6879 -566 6945 -60
rect 7071 -566 7137 -60
rect 7263 -566 7329 -60
rect 7455 -566 7521 -60
rect 7647 -566 7713 -60
rect 7839 -566 7905 -60
rect 8031 -566 8097 -60
rect 8223 -566 8289 -60
rect 8415 -566 8481 -60
rect 8607 -566 8673 -60
rect 8799 -566 8865 -60
rect 8991 -566 9057 -60
rect 9183 -566 9249 -60
rect 9375 -566 9441 -60
rect 9567 -566 9633 -60
rect 9759 -566 9825 -60
rect 9951 -566 10017 -60
rect 10143 -566 10209 -60
rect 10335 -566 10401 -60
rect 10527 -566 10593 -60
<< metal3 >>
rect -10603 -60 -10517 -50
rect -10603 -566 -10593 -60
rect -10527 -566 -10517 -60
rect -10603 -576 -10517 -566
rect -10411 -60 -10325 -50
rect -10411 -566 -10401 -60
rect -10335 -566 -10325 -60
rect -10411 -576 -10325 -566
rect -10219 -60 -10133 -50
rect -10219 -566 -10209 -60
rect -10143 -566 -10133 -60
rect -10219 -576 -10133 -566
rect -10027 -60 -9941 -50
rect -10027 -566 -10017 -60
rect -9951 -566 -9941 -60
rect -10027 -576 -9941 -566
rect -9835 -60 -9749 -50
rect -9835 -566 -9825 -60
rect -9759 -566 -9749 -60
rect -9835 -576 -9749 -566
rect -9643 -60 -9557 -50
rect -9643 -566 -9633 -60
rect -9567 -566 -9557 -60
rect -9643 -576 -9557 -566
rect -9451 -60 -9365 -50
rect -9451 -566 -9441 -60
rect -9375 -566 -9365 -60
rect -9451 -576 -9365 -566
rect -9259 -60 -9173 -50
rect -9259 -566 -9249 -60
rect -9183 -566 -9173 -60
rect -9259 -576 -9173 -566
rect -9067 -60 -8981 -50
rect -9067 -566 -9057 -60
rect -8991 -566 -8981 -60
rect -9067 -576 -8981 -566
rect -8875 -60 -8789 -50
rect -8875 -566 -8865 -60
rect -8799 -566 -8789 -60
rect -8875 -576 -8789 -566
rect -8683 -60 -8597 -50
rect -8683 -566 -8673 -60
rect -8607 -566 -8597 -60
rect -8683 -576 -8597 -566
rect -8491 -60 -8405 -50
rect -8491 -566 -8481 -60
rect -8415 -566 -8405 -60
rect -8491 -576 -8405 -566
rect -8299 -60 -8213 -50
rect -8299 -566 -8289 -60
rect -8223 -566 -8213 -60
rect -8299 -576 -8213 -566
rect -8107 -60 -8021 -50
rect -8107 -566 -8097 -60
rect -8031 -566 -8021 -60
rect -8107 -576 -8021 -566
rect -7915 -60 -7829 -50
rect -7915 -566 -7905 -60
rect -7839 -566 -7829 -60
rect -7915 -576 -7829 -566
rect -7723 -60 -7637 -50
rect -7723 -566 -7713 -60
rect -7647 -566 -7637 -60
rect -7723 -576 -7637 -566
rect -7531 -60 -7445 -50
rect -7531 -566 -7521 -60
rect -7455 -566 -7445 -60
rect -7531 -576 -7445 -566
rect -7339 -60 -7253 -50
rect -7339 -566 -7329 -60
rect -7263 -566 -7253 -60
rect -7339 -576 -7253 -566
rect -7147 -60 -7061 -50
rect -7147 -566 -7137 -60
rect -7071 -566 -7061 -60
rect -7147 -576 -7061 -566
rect -6955 -60 -6869 -50
rect -6955 -566 -6945 -60
rect -6879 -566 -6869 -60
rect -6955 -576 -6869 -566
rect -6763 -60 -6677 -50
rect -6763 -566 -6753 -60
rect -6687 -566 -6677 -60
rect -6763 -576 -6677 -566
rect -6571 -60 -6485 -50
rect -6571 -566 -6561 -60
rect -6495 -566 -6485 -60
rect -6571 -576 -6485 -566
rect -6379 -60 -6293 -50
rect -6379 -566 -6369 -60
rect -6303 -566 -6293 -60
rect -6379 -576 -6293 -566
rect -6187 -60 -6101 -50
rect -6187 -566 -6177 -60
rect -6111 -566 -6101 -60
rect -6187 -576 -6101 -566
rect -5995 -60 -5909 -50
rect -5995 -566 -5985 -60
rect -5919 -566 -5909 -60
rect -5995 -576 -5909 -566
rect -5803 -60 -5717 -50
rect -5803 -566 -5793 -60
rect -5727 -566 -5717 -60
rect -5803 -576 -5717 -566
rect -5611 -60 -5525 -50
rect -5611 -566 -5601 -60
rect -5535 -566 -5525 -60
rect -5611 -576 -5525 -566
rect -5419 -60 -5333 -50
rect -5419 -566 -5409 -60
rect -5343 -566 -5333 -60
rect -5419 -576 -5333 -566
rect -5227 -60 -5141 -50
rect -5227 -566 -5217 -60
rect -5151 -566 -5141 -60
rect -5227 -576 -5141 -566
rect -5035 -60 -4949 -50
rect -5035 -566 -5025 -60
rect -4959 -566 -4949 -60
rect -5035 -576 -4949 -566
rect -4843 -60 -4757 -50
rect -4843 -566 -4833 -60
rect -4767 -566 -4757 -60
rect -4843 -576 -4757 -566
rect -4651 -60 -4565 -50
rect -4651 -566 -4641 -60
rect -4575 -566 -4565 -60
rect -4651 -576 -4565 -566
rect -4459 -60 -4373 -50
rect -4459 -566 -4449 -60
rect -4383 -566 -4373 -60
rect -4459 -576 -4373 -566
rect -4267 -60 -4181 -50
rect -4267 -566 -4257 -60
rect -4191 -566 -4181 -60
rect -4267 -576 -4181 -566
rect -4075 -60 -3989 -50
rect -4075 -566 -4065 -60
rect -3999 -566 -3989 -60
rect -4075 -576 -3989 -566
rect -3883 -60 -3797 -50
rect -3883 -566 -3873 -60
rect -3807 -566 -3797 -60
rect -3883 -576 -3797 -566
rect -3691 -60 -3605 -50
rect -3691 -566 -3681 -60
rect -3615 -566 -3605 -60
rect -3691 -576 -3605 -566
rect -3499 -60 -3413 -50
rect -3499 -566 -3489 -60
rect -3423 -566 -3413 -60
rect -3499 -576 -3413 -566
rect -3307 -60 -3221 -50
rect -3307 -566 -3297 -60
rect -3231 -566 -3221 -60
rect -3307 -576 -3221 -566
rect -3115 -60 -3029 -50
rect -3115 -566 -3105 -60
rect -3039 -566 -3029 -60
rect -3115 -576 -3029 -566
rect -2923 -60 -2837 -50
rect -2923 -566 -2913 -60
rect -2847 -566 -2837 -60
rect -2923 -576 -2837 -566
rect -2731 -60 -2645 -50
rect -2731 -566 -2721 -60
rect -2655 -566 -2645 -60
rect -2731 -576 -2645 -566
rect -2539 -60 -2453 -50
rect -2539 -566 -2529 -60
rect -2463 -566 -2453 -60
rect -2539 -576 -2453 -566
rect -2347 -60 -2261 -50
rect -2347 -566 -2337 -60
rect -2271 -566 -2261 -60
rect -2347 -576 -2261 -566
rect -2155 -60 -2069 -50
rect -2155 -566 -2145 -60
rect -2079 -566 -2069 -60
rect -2155 -576 -2069 -566
rect -1963 -60 -1877 -50
rect -1963 -566 -1953 -60
rect -1887 -566 -1877 -60
rect -1963 -576 -1877 -566
rect -1771 -60 -1685 -50
rect -1771 -566 -1761 -60
rect -1695 -566 -1685 -60
rect -1771 -576 -1685 -566
rect -1579 -60 -1493 -50
rect -1579 -566 -1569 -60
rect -1503 -566 -1493 -60
rect -1579 -576 -1493 -566
rect -1387 -60 -1301 -50
rect -1387 -566 -1377 -60
rect -1311 -566 -1301 -60
rect -1387 -576 -1301 -566
rect -1195 -60 -1109 -50
rect -1195 -566 -1185 -60
rect -1119 -566 -1109 -60
rect -1195 -576 -1109 -566
rect -1003 -60 -917 -50
rect -1003 -566 -993 -60
rect -927 -566 -917 -60
rect -1003 -576 -917 -566
rect -811 -60 -725 -50
rect -811 -566 -801 -60
rect -735 -566 -725 -60
rect -811 -576 -725 -566
rect -619 -60 -533 -50
rect -619 -566 -609 -60
rect -543 -566 -533 -60
rect -619 -576 -533 -566
rect -427 -60 -341 -50
rect -427 -566 -417 -60
rect -351 -566 -341 -60
rect -427 -576 -341 -566
rect -235 -60 -149 -50
rect -235 -566 -225 -60
rect -159 -566 -149 -60
rect -235 -576 -149 -566
rect -43 -60 43 -50
rect -43 -566 -33 -60
rect 33 -566 43 -60
rect -43 -576 43 -566
rect 149 -60 235 -50
rect 149 -566 159 -60
rect 225 -566 235 -60
rect 149 -576 235 -566
rect 341 -60 427 -50
rect 341 -566 351 -60
rect 417 -566 427 -60
rect 341 -576 427 -566
rect 533 -60 619 -50
rect 533 -566 543 -60
rect 609 -566 619 -60
rect 533 -576 619 -566
rect 725 -60 811 -50
rect 725 -566 735 -60
rect 801 -566 811 -60
rect 725 -576 811 -566
rect 917 -60 1003 -50
rect 917 -566 927 -60
rect 993 -566 1003 -60
rect 917 -576 1003 -566
rect 1109 -60 1195 -50
rect 1109 -566 1119 -60
rect 1185 -566 1195 -60
rect 1109 -576 1195 -566
rect 1301 -60 1387 -50
rect 1301 -566 1311 -60
rect 1377 -566 1387 -60
rect 1301 -576 1387 -566
rect 1493 -60 1579 -50
rect 1493 -566 1503 -60
rect 1569 -566 1579 -60
rect 1493 -576 1579 -566
rect 1685 -60 1771 -50
rect 1685 -566 1695 -60
rect 1761 -566 1771 -60
rect 1685 -576 1771 -566
rect 1877 -60 1963 -50
rect 1877 -566 1887 -60
rect 1953 -566 1963 -60
rect 1877 -576 1963 -566
rect 2069 -60 2155 -50
rect 2069 -566 2079 -60
rect 2145 -566 2155 -60
rect 2069 -576 2155 -566
rect 2261 -60 2347 -50
rect 2261 -566 2271 -60
rect 2337 -566 2347 -60
rect 2261 -576 2347 -566
rect 2453 -60 2539 -50
rect 2453 -566 2463 -60
rect 2529 -566 2539 -60
rect 2453 -576 2539 -566
rect 2645 -60 2731 -50
rect 2645 -566 2655 -60
rect 2721 -566 2731 -60
rect 2645 -576 2731 -566
rect 2837 -60 2923 -50
rect 2837 -566 2847 -60
rect 2913 -566 2923 -60
rect 2837 -576 2923 -566
rect 3029 -60 3115 -50
rect 3029 -566 3039 -60
rect 3105 -566 3115 -60
rect 3029 -576 3115 -566
rect 3221 -60 3307 -50
rect 3221 -566 3231 -60
rect 3297 -566 3307 -60
rect 3221 -576 3307 -566
rect 3413 -60 3499 -50
rect 3413 -566 3423 -60
rect 3489 -566 3499 -60
rect 3413 -576 3499 -566
rect 3605 -60 3691 -50
rect 3605 -566 3615 -60
rect 3681 -566 3691 -60
rect 3605 -576 3691 -566
rect 3797 -60 3883 -50
rect 3797 -566 3807 -60
rect 3873 -566 3883 -60
rect 3797 -576 3883 -566
rect 3989 -60 4075 -50
rect 3989 -566 3999 -60
rect 4065 -566 4075 -60
rect 3989 -576 4075 -566
rect 4181 -60 4267 -50
rect 4181 -566 4191 -60
rect 4257 -566 4267 -60
rect 4181 -576 4267 -566
rect 4373 -60 4459 -50
rect 4373 -566 4383 -60
rect 4449 -566 4459 -60
rect 4373 -576 4459 -566
rect 4565 -60 4651 -50
rect 4565 -566 4575 -60
rect 4641 -566 4651 -60
rect 4565 -576 4651 -566
rect 4757 -60 4843 -50
rect 4757 -566 4767 -60
rect 4833 -566 4843 -60
rect 4757 -576 4843 -566
rect 4949 -60 5035 -50
rect 4949 -566 4959 -60
rect 5025 -566 5035 -60
rect 4949 -576 5035 -566
rect 5141 -60 5227 -50
rect 5141 -566 5151 -60
rect 5217 -566 5227 -60
rect 5141 -576 5227 -566
rect 5333 -60 5419 -50
rect 5333 -566 5343 -60
rect 5409 -566 5419 -60
rect 5333 -576 5419 -566
rect 5525 -60 5611 -50
rect 5525 -566 5535 -60
rect 5601 -566 5611 -60
rect 5525 -576 5611 -566
rect 5717 -60 5803 -50
rect 5717 -566 5727 -60
rect 5793 -566 5803 -60
rect 5717 -576 5803 -566
rect 5909 -60 5995 -50
rect 5909 -566 5919 -60
rect 5985 -566 5995 -60
rect 5909 -576 5995 -566
rect 6101 -60 6187 -50
rect 6101 -566 6111 -60
rect 6177 -566 6187 -60
rect 6101 -576 6187 -566
rect 6293 -60 6379 -50
rect 6293 -566 6303 -60
rect 6369 -566 6379 -60
rect 6293 -576 6379 -566
rect 6485 -60 6571 -50
rect 6485 -566 6495 -60
rect 6561 -566 6571 -60
rect 6485 -576 6571 -566
rect 6677 -60 6763 -50
rect 6677 -566 6687 -60
rect 6753 -566 6763 -60
rect 6677 -576 6763 -566
rect 6869 -60 6955 -50
rect 6869 -566 6879 -60
rect 6945 -566 6955 -60
rect 6869 -576 6955 -566
rect 7061 -60 7147 -50
rect 7061 -566 7071 -60
rect 7137 -566 7147 -60
rect 7061 -576 7147 -566
rect 7253 -60 7339 -50
rect 7253 -566 7263 -60
rect 7329 -566 7339 -60
rect 7253 -576 7339 -566
rect 7445 -60 7531 -50
rect 7445 -566 7455 -60
rect 7521 -566 7531 -60
rect 7445 -576 7531 -566
rect 7637 -60 7723 -50
rect 7637 -566 7647 -60
rect 7713 -566 7723 -60
rect 7637 -576 7723 -566
rect 7829 -60 7915 -50
rect 7829 -566 7839 -60
rect 7905 -566 7915 -60
rect 7829 -576 7915 -566
rect 8021 -60 8107 -50
rect 8021 -566 8031 -60
rect 8097 -566 8107 -60
rect 8021 -576 8107 -566
rect 8213 -60 8299 -50
rect 8213 -566 8223 -60
rect 8289 -566 8299 -60
rect 8213 -576 8299 -566
rect 8405 -60 8491 -50
rect 8405 -566 8415 -60
rect 8481 -566 8491 -60
rect 8405 -576 8491 -566
rect 8597 -60 8683 -50
rect 8597 -566 8607 -60
rect 8673 -566 8683 -60
rect 8597 -576 8683 -566
rect 8789 -60 8875 -50
rect 8789 -566 8799 -60
rect 8865 -566 8875 -60
rect 8789 -576 8875 -566
rect 8981 -60 9067 -50
rect 8981 -566 8991 -60
rect 9057 -566 9067 -60
rect 8981 -576 9067 -566
rect 9173 -60 9259 -50
rect 9173 -566 9183 -60
rect 9249 -566 9259 -60
rect 9173 -576 9259 -566
rect 9365 -60 9451 -50
rect 9365 -566 9375 -60
rect 9441 -566 9451 -60
rect 9365 -576 9451 -566
rect 9557 -60 9643 -50
rect 9557 -566 9567 -60
rect 9633 -566 9643 -60
rect 9557 -576 9643 -566
rect 9749 -60 9835 -50
rect 9749 -566 9759 -60
rect 9825 -566 9835 -60
rect 9749 -576 9835 -566
rect 9941 -60 10027 -50
rect 9941 -566 9951 -60
rect 10017 -566 10027 -60
rect 9941 -576 10027 -566
rect 10133 -60 10219 -50
rect 10133 -566 10143 -60
rect 10209 -566 10219 -60
rect 10133 -576 10219 -566
rect 10325 -60 10411 -50
rect 10325 -566 10335 -60
rect 10401 -566 10411 -60
rect 10325 -576 10411 -566
rect 10517 -60 10603 -50
rect 10517 -566 10527 -60
rect 10593 -566 10603 -60
rect 10517 -576 10603 -566
<< via3 >>
rect -10593 -566 -10527 -60
rect -10401 -566 -10335 -60
rect -10209 -566 -10143 -60
rect -10017 -566 -9951 -60
rect -9825 -566 -9759 -60
rect -9633 -566 -9567 -60
rect -9441 -566 -9375 -60
rect -9249 -566 -9183 -60
rect -9057 -566 -8991 -60
rect -8865 -566 -8799 -60
rect -8673 -566 -8607 -60
rect -8481 -566 -8415 -60
rect -8289 -566 -8223 -60
rect -8097 -566 -8031 -60
rect -7905 -566 -7839 -60
rect -7713 -566 -7647 -60
rect -7521 -566 -7455 -60
rect -7329 -566 -7263 -60
rect -7137 -566 -7071 -60
rect -6945 -566 -6879 -60
rect -6753 -566 -6687 -60
rect -6561 -566 -6495 -60
rect -6369 -566 -6303 -60
rect -6177 -566 -6111 -60
rect -5985 -566 -5919 -60
rect -5793 -566 -5727 -60
rect -5601 -566 -5535 -60
rect -5409 -566 -5343 -60
rect -5217 -566 -5151 -60
rect -5025 -566 -4959 -60
rect -4833 -566 -4767 -60
rect -4641 -566 -4575 -60
rect -4449 -566 -4383 -60
rect -4257 -566 -4191 -60
rect -4065 -566 -3999 -60
rect -3873 -566 -3807 -60
rect -3681 -566 -3615 -60
rect -3489 -566 -3423 -60
rect -3297 -566 -3231 -60
rect -3105 -566 -3039 -60
rect -2913 -566 -2847 -60
rect -2721 -566 -2655 -60
rect -2529 -566 -2463 -60
rect -2337 -566 -2271 -60
rect -2145 -566 -2079 -60
rect -1953 -566 -1887 -60
rect -1761 -566 -1695 -60
rect -1569 -566 -1503 -60
rect -1377 -566 -1311 -60
rect -1185 -566 -1119 -60
rect -993 -566 -927 -60
rect -801 -566 -735 -60
rect -609 -566 -543 -60
rect -417 -566 -351 -60
rect -225 -566 -159 -60
rect -33 -566 33 -60
rect 159 -566 225 -60
rect 351 -566 417 -60
rect 543 -566 609 -60
rect 735 -566 801 -60
rect 927 -566 993 -60
rect 1119 -566 1185 -60
rect 1311 -566 1377 -60
rect 1503 -566 1569 -60
rect 1695 -566 1761 -60
rect 1887 -566 1953 -60
rect 2079 -566 2145 -60
rect 2271 -566 2337 -60
rect 2463 -566 2529 -60
rect 2655 -566 2721 -60
rect 2847 -566 2913 -60
rect 3039 -566 3105 -60
rect 3231 -566 3297 -60
rect 3423 -566 3489 -60
rect 3615 -566 3681 -60
rect 3807 -566 3873 -60
rect 3999 -566 4065 -60
rect 4191 -566 4257 -60
rect 4383 -566 4449 -60
rect 4575 -566 4641 -60
rect 4767 -566 4833 -60
rect 4959 -566 5025 -60
rect 5151 -566 5217 -60
rect 5343 -566 5409 -60
rect 5535 -566 5601 -60
rect 5727 -566 5793 -60
rect 5919 -566 5985 -60
rect 6111 -566 6177 -60
rect 6303 -566 6369 -60
rect 6495 -566 6561 -60
rect 6687 -566 6753 -60
rect 6879 -566 6945 -60
rect 7071 -566 7137 -60
rect 7263 -566 7329 -60
rect 7455 -566 7521 -60
rect 7647 -566 7713 -60
rect 7839 -566 7905 -60
rect 8031 -566 8097 -60
rect 8223 -566 8289 -60
rect 8415 -566 8481 -60
rect 8607 -566 8673 -60
rect 8799 -566 8865 -60
rect 8991 -566 9057 -60
rect 9183 -566 9249 -60
rect 9375 -566 9441 -60
rect 9567 -566 9633 -60
rect 9759 -566 9825 -60
rect 9951 -566 10017 -60
rect 10143 -566 10209 -60
rect 10335 -566 10401 -60
rect 10527 -566 10593 -60
<< metal4 >>
rect -10603 -60 -10517 -50
rect -10603 -566 -10593 -60
rect -10527 -566 -10517 -60
rect -10603 -576 -10517 -566
rect -10411 -60 -10325 -50
rect -10411 -566 -10401 -60
rect -10335 -566 -10325 -60
rect -10411 -576 -10325 -566
rect -10219 -60 -10133 -50
rect -10219 -566 -10209 -60
rect -10143 -566 -10133 -60
rect -10219 -576 -10133 -566
rect -10027 -60 -9941 -50
rect -10027 -566 -10017 -60
rect -9951 -566 -9941 -60
rect -10027 -576 -9941 -566
rect -9835 -60 -9749 -50
rect -9835 -566 -9825 -60
rect -9759 -566 -9749 -60
rect -9835 -576 -9749 -566
rect -9643 -60 -9557 -50
rect -9643 -566 -9633 -60
rect -9567 -566 -9557 -60
rect -9643 -576 -9557 -566
rect -9451 -60 -9365 -50
rect -9451 -566 -9441 -60
rect -9375 -566 -9365 -60
rect -9451 -576 -9365 -566
rect -9259 -60 -9173 -50
rect -9259 -566 -9249 -60
rect -9183 -566 -9173 -60
rect -9259 -576 -9173 -566
rect -9067 -60 -8981 -50
rect -9067 -566 -9057 -60
rect -8991 -566 -8981 -60
rect -9067 -576 -8981 -566
rect -8875 -60 -8789 -50
rect -8875 -566 -8865 -60
rect -8799 -566 -8789 -60
rect -8875 -576 -8789 -566
rect -8683 -60 -8597 -50
rect -8683 -566 -8673 -60
rect -8607 -566 -8597 -60
rect -8683 -576 -8597 -566
rect -8491 -60 -8405 -50
rect -8491 -566 -8481 -60
rect -8415 -566 -8405 -60
rect -8491 -576 -8405 -566
rect -8299 -60 -8213 -50
rect -8299 -566 -8289 -60
rect -8223 -566 -8213 -60
rect -8299 -576 -8213 -566
rect -8107 -60 -8021 -50
rect -8107 -566 -8097 -60
rect -8031 -566 -8021 -60
rect -8107 -576 -8021 -566
rect -7915 -60 -7829 -50
rect -7915 -566 -7905 -60
rect -7839 -566 -7829 -60
rect -7915 -576 -7829 -566
rect -7723 -60 -7637 -50
rect -7723 -566 -7713 -60
rect -7647 -566 -7637 -60
rect -7723 -576 -7637 -566
rect -7531 -60 -7445 -50
rect -7531 -566 -7521 -60
rect -7455 -566 -7445 -60
rect -7531 -576 -7445 -566
rect -7339 -60 -7253 -50
rect -7339 -566 -7329 -60
rect -7263 -566 -7253 -60
rect -7339 -576 -7253 -566
rect -7147 -60 -7061 -50
rect -7147 -566 -7137 -60
rect -7071 -566 -7061 -60
rect -7147 -576 -7061 -566
rect -6955 -60 -6869 -50
rect -6955 -566 -6945 -60
rect -6879 -566 -6869 -60
rect -6955 -576 -6869 -566
rect -6763 -60 -6677 -50
rect -6763 -566 -6753 -60
rect -6687 -566 -6677 -60
rect -6763 -576 -6677 -566
rect -6571 -60 -6485 -50
rect -6571 -566 -6561 -60
rect -6495 -566 -6485 -60
rect -6571 -576 -6485 -566
rect -6379 -60 -6293 -50
rect -6379 -566 -6369 -60
rect -6303 -566 -6293 -60
rect -6379 -576 -6293 -566
rect -6187 -60 -6101 -50
rect -6187 -566 -6177 -60
rect -6111 -566 -6101 -60
rect -6187 -576 -6101 -566
rect -5995 -60 -5909 -50
rect -5995 -566 -5985 -60
rect -5919 -566 -5909 -60
rect -5995 -576 -5909 -566
rect -5803 -60 -5717 -50
rect -5803 -566 -5793 -60
rect -5727 -566 -5717 -60
rect -5803 -576 -5717 -566
rect -5611 -60 -5525 -50
rect -5611 -566 -5601 -60
rect -5535 -566 -5525 -60
rect -5611 -576 -5525 -566
rect -5419 -60 -5333 -50
rect -5419 -566 -5409 -60
rect -5343 -566 -5333 -60
rect -5419 -576 -5333 -566
rect -5227 -60 -5141 -50
rect -5227 -566 -5217 -60
rect -5151 -566 -5141 -60
rect -5227 -576 -5141 -566
rect -5035 -60 -4949 -50
rect -5035 -566 -5025 -60
rect -4959 -566 -4949 -60
rect -5035 -576 -4949 -566
rect -4843 -60 -4757 -50
rect -4843 -566 -4833 -60
rect -4767 -566 -4757 -60
rect -4843 -576 -4757 -566
rect -4651 -60 -4565 -50
rect -4651 -566 -4641 -60
rect -4575 -566 -4565 -60
rect -4651 -576 -4565 -566
rect -4459 -60 -4373 -50
rect -4459 -566 -4449 -60
rect -4383 -566 -4373 -60
rect -4459 -576 -4373 -566
rect -4267 -60 -4181 -50
rect -4267 -566 -4257 -60
rect -4191 -566 -4181 -60
rect -4267 -576 -4181 -566
rect -4075 -60 -3989 -50
rect -4075 -566 -4065 -60
rect -3999 -566 -3989 -60
rect -4075 -576 -3989 -566
rect -3883 -60 -3797 -50
rect -3883 -566 -3873 -60
rect -3807 -566 -3797 -60
rect -3883 -576 -3797 -566
rect -3691 -60 -3605 -50
rect -3691 -566 -3681 -60
rect -3615 -566 -3605 -60
rect -3691 -576 -3605 -566
rect -3499 -60 -3413 -50
rect -3499 -566 -3489 -60
rect -3423 -566 -3413 -60
rect -3499 -576 -3413 -566
rect -3307 -60 -3221 -50
rect -3307 -566 -3297 -60
rect -3231 -566 -3221 -60
rect -3307 -576 -3221 -566
rect -3115 -60 -3029 -50
rect -3115 -566 -3105 -60
rect -3039 -566 -3029 -60
rect -3115 -576 -3029 -566
rect -2923 -60 -2837 -50
rect -2923 -566 -2913 -60
rect -2847 -566 -2837 -60
rect -2923 -576 -2837 -566
rect -2731 -60 -2645 -50
rect -2731 -566 -2721 -60
rect -2655 -566 -2645 -60
rect -2731 -576 -2645 -566
rect -2539 -60 -2453 -50
rect -2539 -566 -2529 -60
rect -2463 -566 -2453 -60
rect -2539 -576 -2453 -566
rect -2347 -60 -2261 -50
rect -2347 -566 -2337 -60
rect -2271 -566 -2261 -60
rect -2347 -576 -2261 -566
rect -2155 -60 -2069 -50
rect -2155 -566 -2145 -60
rect -2079 -566 -2069 -60
rect -2155 -576 -2069 -566
rect -1963 -60 -1877 -50
rect -1963 -566 -1953 -60
rect -1887 -566 -1877 -60
rect -1963 -576 -1877 -566
rect -1771 -60 -1685 -50
rect -1771 -566 -1761 -60
rect -1695 -566 -1685 -60
rect -1771 -576 -1685 -566
rect -1579 -60 -1493 -50
rect -1579 -566 -1569 -60
rect -1503 -566 -1493 -60
rect -1579 -576 -1493 -566
rect -1387 -60 -1301 -50
rect -1387 -566 -1377 -60
rect -1311 -566 -1301 -60
rect -1387 -576 -1301 -566
rect -1195 -60 -1109 -50
rect -1195 -566 -1185 -60
rect -1119 -566 -1109 -60
rect -1195 -576 -1109 -566
rect -1003 -60 -917 -50
rect -1003 -566 -993 -60
rect -927 -566 -917 -60
rect -1003 -576 -917 -566
rect -811 -60 -725 -50
rect -811 -566 -801 -60
rect -735 -566 -725 -60
rect -811 -576 -725 -566
rect -619 -60 -533 -50
rect -619 -566 -609 -60
rect -543 -566 -533 -60
rect -619 -576 -533 -566
rect -427 -60 -341 -50
rect -427 -566 -417 -60
rect -351 -566 -341 -60
rect -427 -576 -341 -566
rect -235 -60 -149 -50
rect -235 -566 -225 -60
rect -159 -566 -149 -60
rect -235 -576 -149 -566
rect -43 -60 43 -50
rect -43 -566 -33 -60
rect 33 -566 43 -60
rect -43 -576 43 -566
rect 149 -60 235 -50
rect 149 -566 159 -60
rect 225 -566 235 -60
rect 149 -576 235 -566
rect 341 -60 427 -50
rect 341 -566 351 -60
rect 417 -566 427 -60
rect 341 -576 427 -566
rect 533 -60 619 -50
rect 533 -566 543 -60
rect 609 -566 619 -60
rect 533 -576 619 -566
rect 725 -60 811 -50
rect 725 -566 735 -60
rect 801 -566 811 -60
rect 725 -576 811 -566
rect 917 -60 1003 -50
rect 917 -566 927 -60
rect 993 -566 1003 -60
rect 917 -576 1003 -566
rect 1109 -60 1195 -50
rect 1109 -566 1119 -60
rect 1185 -566 1195 -60
rect 1109 -576 1195 -566
rect 1301 -60 1387 -50
rect 1301 -566 1311 -60
rect 1377 -566 1387 -60
rect 1301 -576 1387 -566
rect 1493 -60 1579 -50
rect 1493 -566 1503 -60
rect 1569 -566 1579 -60
rect 1493 -576 1579 -566
rect 1685 -60 1771 -50
rect 1685 -566 1695 -60
rect 1761 -566 1771 -60
rect 1685 -576 1771 -566
rect 1877 -60 1963 -50
rect 1877 -566 1887 -60
rect 1953 -566 1963 -60
rect 1877 -576 1963 -566
rect 2069 -60 2155 -50
rect 2069 -566 2079 -60
rect 2145 -566 2155 -60
rect 2069 -576 2155 -566
rect 2261 -60 2347 -50
rect 2261 -566 2271 -60
rect 2337 -566 2347 -60
rect 2261 -576 2347 -566
rect 2453 -60 2539 -50
rect 2453 -566 2463 -60
rect 2529 -566 2539 -60
rect 2453 -576 2539 -566
rect 2645 -60 2731 -50
rect 2645 -566 2655 -60
rect 2721 -566 2731 -60
rect 2645 -576 2731 -566
rect 2837 -60 2923 -50
rect 2837 -566 2847 -60
rect 2913 -566 2923 -60
rect 2837 -576 2923 -566
rect 3029 -60 3115 -50
rect 3029 -566 3039 -60
rect 3105 -566 3115 -60
rect 3029 -576 3115 -566
rect 3221 -60 3307 -50
rect 3221 -566 3231 -60
rect 3297 -566 3307 -60
rect 3221 -576 3307 -566
rect 3413 -60 3499 -50
rect 3413 -566 3423 -60
rect 3489 -566 3499 -60
rect 3413 -576 3499 -566
rect 3605 -60 3691 -50
rect 3605 -566 3615 -60
rect 3681 -566 3691 -60
rect 3605 -576 3691 -566
rect 3797 -60 3883 -50
rect 3797 -566 3807 -60
rect 3873 -566 3883 -60
rect 3797 -576 3883 -566
rect 3989 -60 4075 -50
rect 3989 -566 3999 -60
rect 4065 -566 4075 -60
rect 3989 -576 4075 -566
rect 4181 -60 4267 -50
rect 4181 -566 4191 -60
rect 4257 -566 4267 -60
rect 4181 -576 4267 -566
rect 4373 -60 4459 -50
rect 4373 -566 4383 -60
rect 4449 -566 4459 -60
rect 4373 -576 4459 -566
rect 4565 -60 4651 -50
rect 4565 -566 4575 -60
rect 4641 -566 4651 -60
rect 4565 -576 4651 -566
rect 4757 -60 4843 -50
rect 4757 -566 4767 -60
rect 4833 -566 4843 -60
rect 4757 -576 4843 -566
rect 4949 -60 5035 -50
rect 4949 -566 4959 -60
rect 5025 -566 5035 -60
rect 4949 -576 5035 -566
rect 5141 -60 5227 -50
rect 5141 -566 5151 -60
rect 5217 -566 5227 -60
rect 5141 -576 5227 -566
rect 5333 -60 5419 -50
rect 5333 -566 5343 -60
rect 5409 -566 5419 -60
rect 5333 -576 5419 -566
rect 5525 -60 5611 -50
rect 5525 -566 5535 -60
rect 5601 -566 5611 -60
rect 5525 -576 5611 -566
rect 5717 -60 5803 -50
rect 5717 -566 5727 -60
rect 5793 -566 5803 -60
rect 5717 -576 5803 -566
rect 5909 -60 5995 -50
rect 5909 -566 5919 -60
rect 5985 -566 5995 -60
rect 5909 -576 5995 -566
rect 6101 -60 6187 -50
rect 6101 -566 6111 -60
rect 6177 -566 6187 -60
rect 6101 -576 6187 -566
rect 6293 -60 6379 -50
rect 6293 -566 6303 -60
rect 6369 -566 6379 -60
rect 6293 -576 6379 -566
rect 6485 -60 6571 -50
rect 6485 -566 6495 -60
rect 6561 -566 6571 -60
rect 6485 -576 6571 -566
rect 6677 -60 6763 -50
rect 6677 -566 6687 -60
rect 6753 -566 6763 -60
rect 6677 -576 6763 -566
rect 6869 -60 6955 -50
rect 6869 -566 6879 -60
rect 6945 -566 6955 -60
rect 6869 -576 6955 -566
rect 7061 -60 7147 -50
rect 7061 -566 7071 -60
rect 7137 -566 7147 -60
rect 7061 -576 7147 -566
rect 7253 -60 7339 -50
rect 7253 -566 7263 -60
rect 7329 -566 7339 -60
rect 7253 -576 7339 -566
rect 7445 -60 7531 -50
rect 7445 -566 7455 -60
rect 7521 -566 7531 -60
rect 7445 -576 7531 -566
rect 7637 -60 7723 -50
rect 7637 -566 7647 -60
rect 7713 -566 7723 -60
rect 7637 -576 7723 -566
rect 7829 -60 7915 -50
rect 7829 -566 7839 -60
rect 7905 -566 7915 -60
rect 7829 -576 7915 -566
rect 8021 -60 8107 -50
rect 8021 -566 8031 -60
rect 8097 -566 8107 -60
rect 8021 -576 8107 -566
rect 8213 -60 8299 -50
rect 8213 -566 8223 -60
rect 8289 -566 8299 -60
rect 8213 -576 8299 -566
rect 8405 -60 8491 -50
rect 8405 -566 8415 -60
rect 8481 -566 8491 -60
rect 8405 -576 8491 -566
rect 8597 -60 8683 -50
rect 8597 -566 8607 -60
rect 8673 -566 8683 -60
rect 8597 -576 8683 -566
rect 8789 -60 8875 -50
rect 8789 -566 8799 -60
rect 8865 -566 8875 -60
rect 8789 -576 8875 -566
rect 8981 -60 9067 -50
rect 8981 -566 8991 -60
rect 9057 -566 9067 -60
rect 8981 -576 9067 -566
rect 9173 -60 9259 -50
rect 9173 -566 9183 -60
rect 9249 -566 9259 -60
rect 9173 -576 9259 -566
rect 9365 -60 9451 -50
rect 9365 -566 9375 -60
rect 9441 -566 9451 -60
rect 9365 -576 9451 -566
rect 9557 -60 9643 -50
rect 9557 -566 9567 -60
rect 9633 -566 9643 -60
rect 9557 -576 9643 -566
rect 9749 -60 9835 -50
rect 9749 -566 9759 -60
rect 9825 -566 9835 -60
rect 9749 -576 9835 -566
rect 9941 -60 10027 -50
rect 9941 -566 9951 -60
rect 10017 -566 10027 -60
rect 9941 -576 10027 -566
rect 10133 -60 10219 -50
rect 10133 -566 10143 -60
rect 10209 -566 10219 -60
rect 10133 -576 10219 -566
rect 10325 -60 10411 -50
rect 10325 -566 10335 -60
rect 10401 -566 10411 -60
rect 10325 -576 10411 -566
rect 10517 -60 10603 -50
rect 10517 -566 10527 -60
rect 10593 -566 10603 -60
rect 10517 -576 10603 -566
<< properties >>
string FIXED_BBOX -10674 -866 10674 866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 0.15 m 1 nf 220 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
