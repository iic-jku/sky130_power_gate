magic
tech sky130A
magscale 1 2
timestamp 1697193002
<< error_p >>
rect -10445 781 -10387 787
rect -10253 781 -10195 787
rect -10061 781 -10003 787
rect -9869 781 -9811 787
rect -9677 781 -9619 787
rect -9485 781 -9427 787
rect -9293 781 -9235 787
rect -9101 781 -9043 787
rect -8909 781 -8851 787
rect -8717 781 -8659 787
rect -8525 781 -8467 787
rect -8333 781 -8275 787
rect -8141 781 -8083 787
rect -7949 781 -7891 787
rect -7757 781 -7699 787
rect -7565 781 -7507 787
rect -7373 781 -7315 787
rect -7181 781 -7123 787
rect -6989 781 -6931 787
rect -6797 781 -6739 787
rect -6605 781 -6547 787
rect -6413 781 -6355 787
rect -6221 781 -6163 787
rect -6029 781 -5971 787
rect -5837 781 -5779 787
rect -5645 781 -5587 787
rect -5453 781 -5395 787
rect -5261 781 -5203 787
rect -5069 781 -5011 787
rect -4877 781 -4819 787
rect -4685 781 -4627 787
rect -4493 781 -4435 787
rect -4301 781 -4243 787
rect -4109 781 -4051 787
rect -3917 781 -3859 787
rect -3725 781 -3667 787
rect -3533 781 -3475 787
rect -3341 781 -3283 787
rect -3149 781 -3091 787
rect -2957 781 -2899 787
rect -2765 781 -2707 787
rect -2573 781 -2515 787
rect -2381 781 -2323 787
rect -2189 781 -2131 787
rect -1997 781 -1939 787
rect -1805 781 -1747 787
rect -1613 781 -1555 787
rect -1421 781 -1363 787
rect -1229 781 -1171 787
rect -1037 781 -979 787
rect -845 781 -787 787
rect -653 781 -595 787
rect -461 781 -403 787
rect -269 781 -211 787
rect -77 781 -19 787
rect 115 781 173 787
rect 307 781 365 787
rect 499 781 557 787
rect 691 781 749 787
rect 883 781 941 787
rect 1075 781 1133 787
rect 1267 781 1325 787
rect 1459 781 1517 787
rect 1651 781 1709 787
rect 1843 781 1901 787
rect 2035 781 2093 787
rect 2227 781 2285 787
rect 2419 781 2477 787
rect 2611 781 2669 787
rect 2803 781 2861 787
rect 2995 781 3053 787
rect 3187 781 3245 787
rect 3379 781 3437 787
rect 3571 781 3629 787
rect 3763 781 3821 787
rect 3955 781 4013 787
rect 4147 781 4205 787
rect 4339 781 4397 787
rect 4531 781 4589 787
rect 4723 781 4781 787
rect 4915 781 4973 787
rect 5107 781 5165 787
rect 5299 781 5357 787
rect 5491 781 5549 787
rect 5683 781 5741 787
rect 5875 781 5933 787
rect 6067 781 6125 787
rect 6259 781 6317 787
rect 6451 781 6509 787
rect 6643 781 6701 787
rect 6835 781 6893 787
rect 7027 781 7085 787
rect 7219 781 7277 787
rect 7411 781 7469 787
rect 7603 781 7661 787
rect 7795 781 7853 787
rect 7987 781 8045 787
rect 8179 781 8237 787
rect 8371 781 8429 787
rect 8563 781 8621 787
rect 8755 781 8813 787
rect 8947 781 9005 787
rect 9139 781 9197 787
rect 9331 781 9389 787
rect 9523 781 9581 787
rect 9715 781 9773 787
rect 9907 781 9965 787
rect 10099 781 10157 787
rect 10291 781 10349 787
rect 10483 781 10541 787
rect -10445 747 -10433 781
rect -10253 747 -10241 781
rect -10061 747 -10049 781
rect -9869 747 -9857 781
rect -9677 747 -9665 781
rect -9485 747 -9473 781
rect -9293 747 -9281 781
rect -9101 747 -9089 781
rect -8909 747 -8897 781
rect -8717 747 -8705 781
rect -8525 747 -8513 781
rect -8333 747 -8321 781
rect -8141 747 -8129 781
rect -7949 747 -7937 781
rect -7757 747 -7745 781
rect -7565 747 -7553 781
rect -7373 747 -7361 781
rect -7181 747 -7169 781
rect -6989 747 -6977 781
rect -6797 747 -6785 781
rect -6605 747 -6593 781
rect -6413 747 -6401 781
rect -6221 747 -6209 781
rect -6029 747 -6017 781
rect -5837 747 -5825 781
rect -5645 747 -5633 781
rect -5453 747 -5441 781
rect -5261 747 -5249 781
rect -5069 747 -5057 781
rect -4877 747 -4865 781
rect -4685 747 -4673 781
rect -4493 747 -4481 781
rect -4301 747 -4289 781
rect -4109 747 -4097 781
rect -3917 747 -3905 781
rect -3725 747 -3713 781
rect -3533 747 -3521 781
rect -3341 747 -3329 781
rect -3149 747 -3137 781
rect -2957 747 -2945 781
rect -2765 747 -2753 781
rect -2573 747 -2561 781
rect -2381 747 -2369 781
rect -2189 747 -2177 781
rect -1997 747 -1985 781
rect -1805 747 -1793 781
rect -1613 747 -1601 781
rect -1421 747 -1409 781
rect -1229 747 -1217 781
rect -1037 747 -1025 781
rect -845 747 -833 781
rect -653 747 -641 781
rect -461 747 -449 781
rect -269 747 -257 781
rect -77 747 -65 781
rect 115 747 127 781
rect 307 747 319 781
rect 499 747 511 781
rect 691 747 703 781
rect 883 747 895 781
rect 1075 747 1087 781
rect 1267 747 1279 781
rect 1459 747 1471 781
rect 1651 747 1663 781
rect 1843 747 1855 781
rect 2035 747 2047 781
rect 2227 747 2239 781
rect 2419 747 2431 781
rect 2611 747 2623 781
rect 2803 747 2815 781
rect 2995 747 3007 781
rect 3187 747 3199 781
rect 3379 747 3391 781
rect 3571 747 3583 781
rect 3763 747 3775 781
rect 3955 747 3967 781
rect 4147 747 4159 781
rect 4339 747 4351 781
rect 4531 747 4543 781
rect 4723 747 4735 781
rect 4915 747 4927 781
rect 5107 747 5119 781
rect 5299 747 5311 781
rect 5491 747 5503 781
rect 5683 747 5695 781
rect 5875 747 5887 781
rect 6067 747 6079 781
rect 6259 747 6271 781
rect 6451 747 6463 781
rect 6643 747 6655 781
rect 6835 747 6847 781
rect 7027 747 7039 781
rect 7219 747 7231 781
rect 7411 747 7423 781
rect 7603 747 7615 781
rect 7795 747 7807 781
rect 7987 747 7999 781
rect 8179 747 8191 781
rect 8371 747 8383 781
rect 8563 747 8575 781
rect 8755 747 8767 781
rect 8947 747 8959 781
rect 9139 747 9151 781
rect 9331 747 9343 781
rect 9523 747 9535 781
rect 9715 747 9727 781
rect 9907 747 9919 781
rect 10099 747 10111 781
rect 10291 747 10303 781
rect 10483 747 10495 781
rect -10445 741 -10387 747
rect -10253 741 -10195 747
rect -10061 741 -10003 747
rect -9869 741 -9811 747
rect -9677 741 -9619 747
rect -9485 741 -9427 747
rect -9293 741 -9235 747
rect -9101 741 -9043 747
rect -8909 741 -8851 747
rect -8717 741 -8659 747
rect -8525 741 -8467 747
rect -8333 741 -8275 747
rect -8141 741 -8083 747
rect -7949 741 -7891 747
rect -7757 741 -7699 747
rect -7565 741 -7507 747
rect -7373 741 -7315 747
rect -7181 741 -7123 747
rect -6989 741 -6931 747
rect -6797 741 -6739 747
rect -6605 741 -6547 747
rect -6413 741 -6355 747
rect -6221 741 -6163 747
rect -6029 741 -5971 747
rect -5837 741 -5779 747
rect -5645 741 -5587 747
rect -5453 741 -5395 747
rect -5261 741 -5203 747
rect -5069 741 -5011 747
rect -4877 741 -4819 747
rect -4685 741 -4627 747
rect -4493 741 -4435 747
rect -4301 741 -4243 747
rect -4109 741 -4051 747
rect -3917 741 -3859 747
rect -3725 741 -3667 747
rect -3533 741 -3475 747
rect -3341 741 -3283 747
rect -3149 741 -3091 747
rect -2957 741 -2899 747
rect -2765 741 -2707 747
rect -2573 741 -2515 747
rect -2381 741 -2323 747
rect -2189 741 -2131 747
rect -1997 741 -1939 747
rect -1805 741 -1747 747
rect -1613 741 -1555 747
rect -1421 741 -1363 747
rect -1229 741 -1171 747
rect -1037 741 -979 747
rect -845 741 -787 747
rect -653 741 -595 747
rect -461 741 -403 747
rect -269 741 -211 747
rect -77 741 -19 747
rect 115 741 173 747
rect 307 741 365 747
rect 499 741 557 747
rect 691 741 749 747
rect 883 741 941 747
rect 1075 741 1133 747
rect 1267 741 1325 747
rect 1459 741 1517 747
rect 1651 741 1709 747
rect 1843 741 1901 747
rect 2035 741 2093 747
rect 2227 741 2285 747
rect 2419 741 2477 747
rect 2611 741 2669 747
rect 2803 741 2861 747
rect 2995 741 3053 747
rect 3187 741 3245 747
rect 3379 741 3437 747
rect 3571 741 3629 747
rect 3763 741 3821 747
rect 3955 741 4013 747
rect 4147 741 4205 747
rect 4339 741 4397 747
rect 4531 741 4589 747
rect 4723 741 4781 747
rect 4915 741 4973 747
rect 5107 741 5165 747
rect 5299 741 5357 747
rect 5491 741 5549 747
rect 5683 741 5741 747
rect 5875 741 5933 747
rect 6067 741 6125 747
rect 6259 741 6317 747
rect 6451 741 6509 747
rect 6643 741 6701 747
rect 6835 741 6893 747
rect 7027 741 7085 747
rect 7219 741 7277 747
rect 7411 741 7469 747
rect 7603 741 7661 747
rect 7795 741 7853 747
rect 7987 741 8045 747
rect 8179 741 8237 747
rect 8371 741 8429 747
rect 8563 741 8621 747
rect 8755 741 8813 747
rect 8947 741 9005 747
rect 9139 741 9197 747
rect 9331 741 9389 747
rect 9523 741 9581 747
rect 9715 741 9773 747
rect 9907 741 9965 747
rect 10099 741 10157 747
rect 10291 741 10349 747
rect 10483 741 10541 747
rect -10541 -747 -10483 -741
rect -10349 -747 -10291 -741
rect -10157 -747 -10099 -741
rect -9965 -747 -9907 -741
rect -9773 -747 -9715 -741
rect -9581 -747 -9523 -741
rect -9389 -747 -9331 -741
rect -9197 -747 -9139 -741
rect -9005 -747 -8947 -741
rect -8813 -747 -8755 -741
rect -8621 -747 -8563 -741
rect -8429 -747 -8371 -741
rect -8237 -747 -8179 -741
rect -8045 -747 -7987 -741
rect -7853 -747 -7795 -741
rect -7661 -747 -7603 -741
rect -7469 -747 -7411 -741
rect -7277 -747 -7219 -741
rect -7085 -747 -7027 -741
rect -6893 -747 -6835 -741
rect -6701 -747 -6643 -741
rect -6509 -747 -6451 -741
rect -6317 -747 -6259 -741
rect -6125 -747 -6067 -741
rect -5933 -747 -5875 -741
rect -5741 -747 -5683 -741
rect -5549 -747 -5491 -741
rect -5357 -747 -5299 -741
rect -5165 -747 -5107 -741
rect -4973 -747 -4915 -741
rect -4781 -747 -4723 -741
rect -4589 -747 -4531 -741
rect -4397 -747 -4339 -741
rect -4205 -747 -4147 -741
rect -4013 -747 -3955 -741
rect -3821 -747 -3763 -741
rect -3629 -747 -3571 -741
rect -3437 -747 -3379 -741
rect -3245 -747 -3187 -741
rect -3053 -747 -2995 -741
rect -2861 -747 -2803 -741
rect -2669 -747 -2611 -741
rect -2477 -747 -2419 -741
rect -2285 -747 -2227 -741
rect -2093 -747 -2035 -741
rect -1901 -747 -1843 -741
rect -1709 -747 -1651 -741
rect -1517 -747 -1459 -741
rect -1325 -747 -1267 -741
rect -1133 -747 -1075 -741
rect -941 -747 -883 -741
rect -749 -747 -691 -741
rect -557 -747 -499 -741
rect -365 -747 -307 -741
rect -173 -747 -115 -741
rect 19 -747 77 -741
rect 211 -747 269 -741
rect 403 -747 461 -741
rect 595 -747 653 -741
rect 787 -747 845 -741
rect 979 -747 1037 -741
rect 1171 -747 1229 -741
rect 1363 -747 1421 -741
rect 1555 -747 1613 -741
rect 1747 -747 1805 -741
rect 1939 -747 1997 -741
rect 2131 -747 2189 -741
rect 2323 -747 2381 -741
rect 2515 -747 2573 -741
rect 2707 -747 2765 -741
rect 2899 -747 2957 -741
rect 3091 -747 3149 -741
rect 3283 -747 3341 -741
rect 3475 -747 3533 -741
rect 3667 -747 3725 -741
rect 3859 -747 3917 -741
rect 4051 -747 4109 -741
rect 4243 -747 4301 -741
rect 4435 -747 4493 -741
rect 4627 -747 4685 -741
rect 4819 -747 4877 -741
rect 5011 -747 5069 -741
rect 5203 -747 5261 -741
rect 5395 -747 5453 -741
rect 5587 -747 5645 -741
rect 5779 -747 5837 -741
rect 5971 -747 6029 -741
rect 6163 -747 6221 -741
rect 6355 -747 6413 -741
rect 6547 -747 6605 -741
rect 6739 -747 6797 -741
rect 6931 -747 6989 -741
rect 7123 -747 7181 -741
rect 7315 -747 7373 -741
rect 7507 -747 7565 -741
rect 7699 -747 7757 -741
rect 7891 -747 7949 -741
rect 8083 -747 8141 -741
rect 8275 -747 8333 -741
rect 8467 -747 8525 -741
rect 8659 -747 8717 -741
rect 8851 -747 8909 -741
rect 9043 -747 9101 -741
rect 9235 -747 9293 -741
rect 9427 -747 9485 -741
rect 9619 -747 9677 -741
rect 9811 -747 9869 -741
rect 10003 -747 10061 -741
rect 10195 -747 10253 -741
rect 10387 -747 10445 -741
rect -10541 -781 -10529 -747
rect -10349 -781 -10337 -747
rect -10157 -781 -10145 -747
rect -9965 -781 -9953 -747
rect -9773 -781 -9761 -747
rect -9581 -781 -9569 -747
rect -9389 -781 -9377 -747
rect -9197 -781 -9185 -747
rect -9005 -781 -8993 -747
rect -8813 -781 -8801 -747
rect -8621 -781 -8609 -747
rect -8429 -781 -8417 -747
rect -8237 -781 -8225 -747
rect -8045 -781 -8033 -747
rect -7853 -781 -7841 -747
rect -7661 -781 -7649 -747
rect -7469 -781 -7457 -747
rect -7277 -781 -7265 -747
rect -7085 -781 -7073 -747
rect -6893 -781 -6881 -747
rect -6701 -781 -6689 -747
rect -6509 -781 -6497 -747
rect -6317 -781 -6305 -747
rect -6125 -781 -6113 -747
rect -5933 -781 -5921 -747
rect -5741 -781 -5729 -747
rect -5549 -781 -5537 -747
rect -5357 -781 -5345 -747
rect -5165 -781 -5153 -747
rect -4973 -781 -4961 -747
rect -4781 -781 -4769 -747
rect -4589 -781 -4577 -747
rect -4397 -781 -4385 -747
rect -4205 -781 -4193 -747
rect -4013 -781 -4001 -747
rect -3821 -781 -3809 -747
rect -3629 -781 -3617 -747
rect -3437 -781 -3425 -747
rect -3245 -781 -3233 -747
rect -3053 -781 -3041 -747
rect -2861 -781 -2849 -747
rect -2669 -781 -2657 -747
rect -2477 -781 -2465 -747
rect -2285 -781 -2273 -747
rect -2093 -781 -2081 -747
rect -1901 -781 -1889 -747
rect -1709 -781 -1697 -747
rect -1517 -781 -1505 -747
rect -1325 -781 -1313 -747
rect -1133 -781 -1121 -747
rect -941 -781 -929 -747
rect -749 -781 -737 -747
rect -557 -781 -545 -747
rect -365 -781 -353 -747
rect -173 -781 -161 -747
rect 19 -781 31 -747
rect 211 -781 223 -747
rect 403 -781 415 -747
rect 595 -781 607 -747
rect 787 -781 799 -747
rect 979 -781 991 -747
rect 1171 -781 1183 -747
rect 1363 -781 1375 -747
rect 1555 -781 1567 -747
rect 1747 -781 1759 -747
rect 1939 -781 1951 -747
rect 2131 -781 2143 -747
rect 2323 -781 2335 -747
rect 2515 -781 2527 -747
rect 2707 -781 2719 -747
rect 2899 -781 2911 -747
rect 3091 -781 3103 -747
rect 3283 -781 3295 -747
rect 3475 -781 3487 -747
rect 3667 -781 3679 -747
rect 3859 -781 3871 -747
rect 4051 -781 4063 -747
rect 4243 -781 4255 -747
rect 4435 -781 4447 -747
rect 4627 -781 4639 -747
rect 4819 -781 4831 -747
rect 5011 -781 5023 -747
rect 5203 -781 5215 -747
rect 5395 -781 5407 -747
rect 5587 -781 5599 -747
rect 5779 -781 5791 -747
rect 5971 -781 5983 -747
rect 6163 -781 6175 -747
rect 6355 -781 6367 -747
rect 6547 -781 6559 -747
rect 6739 -781 6751 -747
rect 6931 -781 6943 -747
rect 7123 -781 7135 -747
rect 7315 -781 7327 -747
rect 7507 -781 7519 -747
rect 7699 -781 7711 -747
rect 7891 -781 7903 -747
rect 8083 -781 8095 -747
rect 8275 -781 8287 -747
rect 8467 -781 8479 -747
rect 8659 -781 8671 -747
rect 8851 -781 8863 -747
rect 9043 -781 9055 -747
rect 9235 -781 9247 -747
rect 9427 -781 9439 -747
rect 9619 -781 9631 -747
rect 9811 -781 9823 -747
rect 10003 -781 10015 -747
rect 10195 -781 10207 -747
rect 10387 -781 10399 -747
rect -10541 -787 -10483 -781
rect -10349 -787 -10291 -781
rect -10157 -787 -10099 -781
rect -9965 -787 -9907 -781
rect -9773 -787 -9715 -781
rect -9581 -787 -9523 -781
rect -9389 -787 -9331 -781
rect -9197 -787 -9139 -781
rect -9005 -787 -8947 -781
rect -8813 -787 -8755 -781
rect -8621 -787 -8563 -781
rect -8429 -787 -8371 -781
rect -8237 -787 -8179 -781
rect -8045 -787 -7987 -781
rect -7853 -787 -7795 -781
rect -7661 -787 -7603 -781
rect -7469 -787 -7411 -781
rect -7277 -787 -7219 -781
rect -7085 -787 -7027 -781
rect -6893 -787 -6835 -781
rect -6701 -787 -6643 -781
rect -6509 -787 -6451 -781
rect -6317 -787 -6259 -781
rect -6125 -787 -6067 -781
rect -5933 -787 -5875 -781
rect -5741 -787 -5683 -781
rect -5549 -787 -5491 -781
rect -5357 -787 -5299 -781
rect -5165 -787 -5107 -781
rect -4973 -787 -4915 -781
rect -4781 -787 -4723 -781
rect -4589 -787 -4531 -781
rect -4397 -787 -4339 -781
rect -4205 -787 -4147 -781
rect -4013 -787 -3955 -781
rect -3821 -787 -3763 -781
rect -3629 -787 -3571 -781
rect -3437 -787 -3379 -781
rect -3245 -787 -3187 -781
rect -3053 -787 -2995 -781
rect -2861 -787 -2803 -781
rect -2669 -787 -2611 -781
rect -2477 -787 -2419 -781
rect -2285 -787 -2227 -781
rect -2093 -787 -2035 -781
rect -1901 -787 -1843 -781
rect -1709 -787 -1651 -781
rect -1517 -787 -1459 -781
rect -1325 -787 -1267 -781
rect -1133 -787 -1075 -781
rect -941 -787 -883 -781
rect -749 -787 -691 -781
rect -557 -787 -499 -781
rect -365 -787 -307 -781
rect -173 -787 -115 -781
rect 19 -787 77 -781
rect 211 -787 269 -781
rect 403 -787 461 -781
rect 595 -787 653 -781
rect 787 -787 845 -781
rect 979 -787 1037 -781
rect 1171 -787 1229 -781
rect 1363 -787 1421 -781
rect 1555 -787 1613 -781
rect 1747 -787 1805 -781
rect 1939 -787 1997 -781
rect 2131 -787 2189 -781
rect 2323 -787 2381 -781
rect 2515 -787 2573 -781
rect 2707 -787 2765 -781
rect 2899 -787 2957 -781
rect 3091 -787 3149 -781
rect 3283 -787 3341 -781
rect 3475 -787 3533 -781
rect 3667 -787 3725 -781
rect 3859 -787 3917 -781
rect 4051 -787 4109 -781
rect 4243 -787 4301 -781
rect 4435 -787 4493 -781
rect 4627 -787 4685 -781
rect 4819 -787 4877 -781
rect 5011 -787 5069 -781
rect 5203 -787 5261 -781
rect 5395 -787 5453 -781
rect 5587 -787 5645 -781
rect 5779 -787 5837 -781
rect 5971 -787 6029 -781
rect 6163 -787 6221 -781
rect 6355 -787 6413 -781
rect 6547 -787 6605 -781
rect 6739 -787 6797 -781
rect 6931 -787 6989 -781
rect 7123 -787 7181 -781
rect 7315 -787 7373 -781
rect 7507 -787 7565 -781
rect 7699 -787 7757 -781
rect 7891 -787 7949 -781
rect 8083 -787 8141 -781
rect 8275 -787 8333 -781
rect 8467 -787 8525 -781
rect 8659 -787 8717 -781
rect 8851 -787 8909 -781
rect 9043 -787 9101 -781
rect 9235 -787 9293 -781
rect 9427 -787 9485 -781
rect 9619 -787 9677 -781
rect 9811 -787 9869 -781
rect 10003 -787 10061 -781
rect 10195 -787 10253 -781
rect 10387 -787 10445 -781
<< nwell >>
rect -10727 -919 10727 919
<< pmos >>
rect -10527 -700 -10497 700
rect -10431 -700 -10401 700
rect -10335 -700 -10305 700
rect -10239 -700 -10209 700
rect -10143 -700 -10113 700
rect -10047 -700 -10017 700
rect -9951 -700 -9921 700
rect -9855 -700 -9825 700
rect -9759 -700 -9729 700
rect -9663 -700 -9633 700
rect -9567 -700 -9537 700
rect -9471 -700 -9441 700
rect -9375 -700 -9345 700
rect -9279 -700 -9249 700
rect -9183 -700 -9153 700
rect -9087 -700 -9057 700
rect -8991 -700 -8961 700
rect -8895 -700 -8865 700
rect -8799 -700 -8769 700
rect -8703 -700 -8673 700
rect -8607 -700 -8577 700
rect -8511 -700 -8481 700
rect -8415 -700 -8385 700
rect -8319 -700 -8289 700
rect -8223 -700 -8193 700
rect -8127 -700 -8097 700
rect -8031 -700 -8001 700
rect -7935 -700 -7905 700
rect -7839 -700 -7809 700
rect -7743 -700 -7713 700
rect -7647 -700 -7617 700
rect -7551 -700 -7521 700
rect -7455 -700 -7425 700
rect -7359 -700 -7329 700
rect -7263 -700 -7233 700
rect -7167 -700 -7137 700
rect -7071 -700 -7041 700
rect -6975 -700 -6945 700
rect -6879 -700 -6849 700
rect -6783 -700 -6753 700
rect -6687 -700 -6657 700
rect -6591 -700 -6561 700
rect -6495 -700 -6465 700
rect -6399 -700 -6369 700
rect -6303 -700 -6273 700
rect -6207 -700 -6177 700
rect -6111 -700 -6081 700
rect -6015 -700 -5985 700
rect -5919 -700 -5889 700
rect -5823 -700 -5793 700
rect -5727 -700 -5697 700
rect -5631 -700 -5601 700
rect -5535 -700 -5505 700
rect -5439 -700 -5409 700
rect -5343 -700 -5313 700
rect -5247 -700 -5217 700
rect -5151 -700 -5121 700
rect -5055 -700 -5025 700
rect -4959 -700 -4929 700
rect -4863 -700 -4833 700
rect -4767 -700 -4737 700
rect -4671 -700 -4641 700
rect -4575 -700 -4545 700
rect -4479 -700 -4449 700
rect -4383 -700 -4353 700
rect -4287 -700 -4257 700
rect -4191 -700 -4161 700
rect -4095 -700 -4065 700
rect -3999 -700 -3969 700
rect -3903 -700 -3873 700
rect -3807 -700 -3777 700
rect -3711 -700 -3681 700
rect -3615 -700 -3585 700
rect -3519 -700 -3489 700
rect -3423 -700 -3393 700
rect -3327 -700 -3297 700
rect -3231 -700 -3201 700
rect -3135 -700 -3105 700
rect -3039 -700 -3009 700
rect -2943 -700 -2913 700
rect -2847 -700 -2817 700
rect -2751 -700 -2721 700
rect -2655 -700 -2625 700
rect -2559 -700 -2529 700
rect -2463 -700 -2433 700
rect -2367 -700 -2337 700
rect -2271 -700 -2241 700
rect -2175 -700 -2145 700
rect -2079 -700 -2049 700
rect -1983 -700 -1953 700
rect -1887 -700 -1857 700
rect -1791 -700 -1761 700
rect -1695 -700 -1665 700
rect -1599 -700 -1569 700
rect -1503 -700 -1473 700
rect -1407 -700 -1377 700
rect -1311 -700 -1281 700
rect -1215 -700 -1185 700
rect -1119 -700 -1089 700
rect -1023 -700 -993 700
rect -927 -700 -897 700
rect -831 -700 -801 700
rect -735 -700 -705 700
rect -639 -700 -609 700
rect -543 -700 -513 700
rect -447 -700 -417 700
rect -351 -700 -321 700
rect -255 -700 -225 700
rect -159 -700 -129 700
rect -63 -700 -33 700
rect 33 -700 63 700
rect 129 -700 159 700
rect 225 -700 255 700
rect 321 -700 351 700
rect 417 -700 447 700
rect 513 -700 543 700
rect 609 -700 639 700
rect 705 -700 735 700
rect 801 -700 831 700
rect 897 -700 927 700
rect 993 -700 1023 700
rect 1089 -700 1119 700
rect 1185 -700 1215 700
rect 1281 -700 1311 700
rect 1377 -700 1407 700
rect 1473 -700 1503 700
rect 1569 -700 1599 700
rect 1665 -700 1695 700
rect 1761 -700 1791 700
rect 1857 -700 1887 700
rect 1953 -700 1983 700
rect 2049 -700 2079 700
rect 2145 -700 2175 700
rect 2241 -700 2271 700
rect 2337 -700 2367 700
rect 2433 -700 2463 700
rect 2529 -700 2559 700
rect 2625 -700 2655 700
rect 2721 -700 2751 700
rect 2817 -700 2847 700
rect 2913 -700 2943 700
rect 3009 -700 3039 700
rect 3105 -700 3135 700
rect 3201 -700 3231 700
rect 3297 -700 3327 700
rect 3393 -700 3423 700
rect 3489 -700 3519 700
rect 3585 -700 3615 700
rect 3681 -700 3711 700
rect 3777 -700 3807 700
rect 3873 -700 3903 700
rect 3969 -700 3999 700
rect 4065 -700 4095 700
rect 4161 -700 4191 700
rect 4257 -700 4287 700
rect 4353 -700 4383 700
rect 4449 -700 4479 700
rect 4545 -700 4575 700
rect 4641 -700 4671 700
rect 4737 -700 4767 700
rect 4833 -700 4863 700
rect 4929 -700 4959 700
rect 5025 -700 5055 700
rect 5121 -700 5151 700
rect 5217 -700 5247 700
rect 5313 -700 5343 700
rect 5409 -700 5439 700
rect 5505 -700 5535 700
rect 5601 -700 5631 700
rect 5697 -700 5727 700
rect 5793 -700 5823 700
rect 5889 -700 5919 700
rect 5985 -700 6015 700
rect 6081 -700 6111 700
rect 6177 -700 6207 700
rect 6273 -700 6303 700
rect 6369 -700 6399 700
rect 6465 -700 6495 700
rect 6561 -700 6591 700
rect 6657 -700 6687 700
rect 6753 -700 6783 700
rect 6849 -700 6879 700
rect 6945 -700 6975 700
rect 7041 -700 7071 700
rect 7137 -700 7167 700
rect 7233 -700 7263 700
rect 7329 -700 7359 700
rect 7425 -700 7455 700
rect 7521 -700 7551 700
rect 7617 -700 7647 700
rect 7713 -700 7743 700
rect 7809 -700 7839 700
rect 7905 -700 7935 700
rect 8001 -700 8031 700
rect 8097 -700 8127 700
rect 8193 -700 8223 700
rect 8289 -700 8319 700
rect 8385 -700 8415 700
rect 8481 -700 8511 700
rect 8577 -700 8607 700
rect 8673 -700 8703 700
rect 8769 -700 8799 700
rect 8865 -700 8895 700
rect 8961 -700 8991 700
rect 9057 -700 9087 700
rect 9153 -700 9183 700
rect 9249 -700 9279 700
rect 9345 -700 9375 700
rect 9441 -700 9471 700
rect 9537 -700 9567 700
rect 9633 -700 9663 700
rect 9729 -700 9759 700
rect 9825 -700 9855 700
rect 9921 -700 9951 700
rect 10017 -700 10047 700
rect 10113 -700 10143 700
rect 10209 -700 10239 700
rect 10305 -700 10335 700
rect 10401 -700 10431 700
rect 10497 -700 10527 700
<< pdiff >>
rect -10589 688 -10527 700
rect -10589 -688 -10577 688
rect -10543 -688 -10527 688
rect -10589 -700 -10527 -688
rect -10497 688 -10431 700
rect -10497 -688 -10481 688
rect -10447 -688 -10431 688
rect -10497 -700 -10431 -688
rect -10401 688 -10335 700
rect -10401 -688 -10385 688
rect -10351 -688 -10335 688
rect -10401 -700 -10335 -688
rect -10305 688 -10239 700
rect -10305 -688 -10289 688
rect -10255 -688 -10239 688
rect -10305 -700 -10239 -688
rect -10209 688 -10143 700
rect -10209 -688 -10193 688
rect -10159 -688 -10143 688
rect -10209 -700 -10143 -688
rect -10113 688 -10047 700
rect -10113 -688 -10097 688
rect -10063 -688 -10047 688
rect -10113 -700 -10047 -688
rect -10017 688 -9951 700
rect -10017 -688 -10001 688
rect -9967 -688 -9951 688
rect -10017 -700 -9951 -688
rect -9921 688 -9855 700
rect -9921 -688 -9905 688
rect -9871 -688 -9855 688
rect -9921 -700 -9855 -688
rect -9825 688 -9759 700
rect -9825 -688 -9809 688
rect -9775 -688 -9759 688
rect -9825 -700 -9759 -688
rect -9729 688 -9663 700
rect -9729 -688 -9713 688
rect -9679 -688 -9663 688
rect -9729 -700 -9663 -688
rect -9633 688 -9567 700
rect -9633 -688 -9617 688
rect -9583 -688 -9567 688
rect -9633 -700 -9567 -688
rect -9537 688 -9471 700
rect -9537 -688 -9521 688
rect -9487 -688 -9471 688
rect -9537 -700 -9471 -688
rect -9441 688 -9375 700
rect -9441 -688 -9425 688
rect -9391 -688 -9375 688
rect -9441 -700 -9375 -688
rect -9345 688 -9279 700
rect -9345 -688 -9329 688
rect -9295 -688 -9279 688
rect -9345 -700 -9279 -688
rect -9249 688 -9183 700
rect -9249 -688 -9233 688
rect -9199 -688 -9183 688
rect -9249 -700 -9183 -688
rect -9153 688 -9087 700
rect -9153 -688 -9137 688
rect -9103 -688 -9087 688
rect -9153 -700 -9087 -688
rect -9057 688 -8991 700
rect -9057 -688 -9041 688
rect -9007 -688 -8991 688
rect -9057 -700 -8991 -688
rect -8961 688 -8895 700
rect -8961 -688 -8945 688
rect -8911 -688 -8895 688
rect -8961 -700 -8895 -688
rect -8865 688 -8799 700
rect -8865 -688 -8849 688
rect -8815 -688 -8799 688
rect -8865 -700 -8799 -688
rect -8769 688 -8703 700
rect -8769 -688 -8753 688
rect -8719 -688 -8703 688
rect -8769 -700 -8703 -688
rect -8673 688 -8607 700
rect -8673 -688 -8657 688
rect -8623 -688 -8607 688
rect -8673 -700 -8607 -688
rect -8577 688 -8511 700
rect -8577 -688 -8561 688
rect -8527 -688 -8511 688
rect -8577 -700 -8511 -688
rect -8481 688 -8415 700
rect -8481 -688 -8465 688
rect -8431 -688 -8415 688
rect -8481 -700 -8415 -688
rect -8385 688 -8319 700
rect -8385 -688 -8369 688
rect -8335 -688 -8319 688
rect -8385 -700 -8319 -688
rect -8289 688 -8223 700
rect -8289 -688 -8273 688
rect -8239 -688 -8223 688
rect -8289 -700 -8223 -688
rect -8193 688 -8127 700
rect -8193 -688 -8177 688
rect -8143 -688 -8127 688
rect -8193 -700 -8127 -688
rect -8097 688 -8031 700
rect -8097 -688 -8081 688
rect -8047 -688 -8031 688
rect -8097 -700 -8031 -688
rect -8001 688 -7935 700
rect -8001 -688 -7985 688
rect -7951 -688 -7935 688
rect -8001 -700 -7935 -688
rect -7905 688 -7839 700
rect -7905 -688 -7889 688
rect -7855 -688 -7839 688
rect -7905 -700 -7839 -688
rect -7809 688 -7743 700
rect -7809 -688 -7793 688
rect -7759 -688 -7743 688
rect -7809 -700 -7743 -688
rect -7713 688 -7647 700
rect -7713 -688 -7697 688
rect -7663 -688 -7647 688
rect -7713 -700 -7647 -688
rect -7617 688 -7551 700
rect -7617 -688 -7601 688
rect -7567 -688 -7551 688
rect -7617 -700 -7551 -688
rect -7521 688 -7455 700
rect -7521 -688 -7505 688
rect -7471 -688 -7455 688
rect -7521 -700 -7455 -688
rect -7425 688 -7359 700
rect -7425 -688 -7409 688
rect -7375 -688 -7359 688
rect -7425 -700 -7359 -688
rect -7329 688 -7263 700
rect -7329 -688 -7313 688
rect -7279 -688 -7263 688
rect -7329 -700 -7263 -688
rect -7233 688 -7167 700
rect -7233 -688 -7217 688
rect -7183 -688 -7167 688
rect -7233 -700 -7167 -688
rect -7137 688 -7071 700
rect -7137 -688 -7121 688
rect -7087 -688 -7071 688
rect -7137 -700 -7071 -688
rect -7041 688 -6975 700
rect -7041 -688 -7025 688
rect -6991 -688 -6975 688
rect -7041 -700 -6975 -688
rect -6945 688 -6879 700
rect -6945 -688 -6929 688
rect -6895 -688 -6879 688
rect -6945 -700 -6879 -688
rect -6849 688 -6783 700
rect -6849 -688 -6833 688
rect -6799 -688 -6783 688
rect -6849 -700 -6783 -688
rect -6753 688 -6687 700
rect -6753 -688 -6737 688
rect -6703 -688 -6687 688
rect -6753 -700 -6687 -688
rect -6657 688 -6591 700
rect -6657 -688 -6641 688
rect -6607 -688 -6591 688
rect -6657 -700 -6591 -688
rect -6561 688 -6495 700
rect -6561 -688 -6545 688
rect -6511 -688 -6495 688
rect -6561 -700 -6495 -688
rect -6465 688 -6399 700
rect -6465 -688 -6449 688
rect -6415 -688 -6399 688
rect -6465 -700 -6399 -688
rect -6369 688 -6303 700
rect -6369 -688 -6353 688
rect -6319 -688 -6303 688
rect -6369 -700 -6303 -688
rect -6273 688 -6207 700
rect -6273 -688 -6257 688
rect -6223 -688 -6207 688
rect -6273 -700 -6207 -688
rect -6177 688 -6111 700
rect -6177 -688 -6161 688
rect -6127 -688 -6111 688
rect -6177 -700 -6111 -688
rect -6081 688 -6015 700
rect -6081 -688 -6065 688
rect -6031 -688 -6015 688
rect -6081 -700 -6015 -688
rect -5985 688 -5919 700
rect -5985 -688 -5969 688
rect -5935 -688 -5919 688
rect -5985 -700 -5919 -688
rect -5889 688 -5823 700
rect -5889 -688 -5873 688
rect -5839 -688 -5823 688
rect -5889 -700 -5823 -688
rect -5793 688 -5727 700
rect -5793 -688 -5777 688
rect -5743 -688 -5727 688
rect -5793 -700 -5727 -688
rect -5697 688 -5631 700
rect -5697 -688 -5681 688
rect -5647 -688 -5631 688
rect -5697 -700 -5631 -688
rect -5601 688 -5535 700
rect -5601 -688 -5585 688
rect -5551 -688 -5535 688
rect -5601 -700 -5535 -688
rect -5505 688 -5439 700
rect -5505 -688 -5489 688
rect -5455 -688 -5439 688
rect -5505 -700 -5439 -688
rect -5409 688 -5343 700
rect -5409 -688 -5393 688
rect -5359 -688 -5343 688
rect -5409 -700 -5343 -688
rect -5313 688 -5247 700
rect -5313 -688 -5297 688
rect -5263 -688 -5247 688
rect -5313 -700 -5247 -688
rect -5217 688 -5151 700
rect -5217 -688 -5201 688
rect -5167 -688 -5151 688
rect -5217 -700 -5151 -688
rect -5121 688 -5055 700
rect -5121 -688 -5105 688
rect -5071 -688 -5055 688
rect -5121 -700 -5055 -688
rect -5025 688 -4959 700
rect -5025 -688 -5009 688
rect -4975 -688 -4959 688
rect -5025 -700 -4959 -688
rect -4929 688 -4863 700
rect -4929 -688 -4913 688
rect -4879 -688 -4863 688
rect -4929 -700 -4863 -688
rect -4833 688 -4767 700
rect -4833 -688 -4817 688
rect -4783 -688 -4767 688
rect -4833 -700 -4767 -688
rect -4737 688 -4671 700
rect -4737 -688 -4721 688
rect -4687 -688 -4671 688
rect -4737 -700 -4671 -688
rect -4641 688 -4575 700
rect -4641 -688 -4625 688
rect -4591 -688 -4575 688
rect -4641 -700 -4575 -688
rect -4545 688 -4479 700
rect -4545 -688 -4529 688
rect -4495 -688 -4479 688
rect -4545 -700 -4479 -688
rect -4449 688 -4383 700
rect -4449 -688 -4433 688
rect -4399 -688 -4383 688
rect -4449 -700 -4383 -688
rect -4353 688 -4287 700
rect -4353 -688 -4337 688
rect -4303 -688 -4287 688
rect -4353 -700 -4287 -688
rect -4257 688 -4191 700
rect -4257 -688 -4241 688
rect -4207 -688 -4191 688
rect -4257 -700 -4191 -688
rect -4161 688 -4095 700
rect -4161 -688 -4145 688
rect -4111 -688 -4095 688
rect -4161 -700 -4095 -688
rect -4065 688 -3999 700
rect -4065 -688 -4049 688
rect -4015 -688 -3999 688
rect -4065 -700 -3999 -688
rect -3969 688 -3903 700
rect -3969 -688 -3953 688
rect -3919 -688 -3903 688
rect -3969 -700 -3903 -688
rect -3873 688 -3807 700
rect -3873 -688 -3857 688
rect -3823 -688 -3807 688
rect -3873 -700 -3807 -688
rect -3777 688 -3711 700
rect -3777 -688 -3761 688
rect -3727 -688 -3711 688
rect -3777 -700 -3711 -688
rect -3681 688 -3615 700
rect -3681 -688 -3665 688
rect -3631 -688 -3615 688
rect -3681 -700 -3615 -688
rect -3585 688 -3519 700
rect -3585 -688 -3569 688
rect -3535 -688 -3519 688
rect -3585 -700 -3519 -688
rect -3489 688 -3423 700
rect -3489 -688 -3473 688
rect -3439 -688 -3423 688
rect -3489 -700 -3423 -688
rect -3393 688 -3327 700
rect -3393 -688 -3377 688
rect -3343 -688 -3327 688
rect -3393 -700 -3327 -688
rect -3297 688 -3231 700
rect -3297 -688 -3281 688
rect -3247 -688 -3231 688
rect -3297 -700 -3231 -688
rect -3201 688 -3135 700
rect -3201 -688 -3185 688
rect -3151 -688 -3135 688
rect -3201 -700 -3135 -688
rect -3105 688 -3039 700
rect -3105 -688 -3089 688
rect -3055 -688 -3039 688
rect -3105 -700 -3039 -688
rect -3009 688 -2943 700
rect -3009 -688 -2993 688
rect -2959 -688 -2943 688
rect -3009 -700 -2943 -688
rect -2913 688 -2847 700
rect -2913 -688 -2897 688
rect -2863 -688 -2847 688
rect -2913 -700 -2847 -688
rect -2817 688 -2751 700
rect -2817 -688 -2801 688
rect -2767 -688 -2751 688
rect -2817 -700 -2751 -688
rect -2721 688 -2655 700
rect -2721 -688 -2705 688
rect -2671 -688 -2655 688
rect -2721 -700 -2655 -688
rect -2625 688 -2559 700
rect -2625 -688 -2609 688
rect -2575 -688 -2559 688
rect -2625 -700 -2559 -688
rect -2529 688 -2463 700
rect -2529 -688 -2513 688
rect -2479 -688 -2463 688
rect -2529 -700 -2463 -688
rect -2433 688 -2367 700
rect -2433 -688 -2417 688
rect -2383 -688 -2367 688
rect -2433 -700 -2367 -688
rect -2337 688 -2271 700
rect -2337 -688 -2321 688
rect -2287 -688 -2271 688
rect -2337 -700 -2271 -688
rect -2241 688 -2175 700
rect -2241 -688 -2225 688
rect -2191 -688 -2175 688
rect -2241 -700 -2175 -688
rect -2145 688 -2079 700
rect -2145 -688 -2129 688
rect -2095 -688 -2079 688
rect -2145 -700 -2079 -688
rect -2049 688 -1983 700
rect -2049 -688 -2033 688
rect -1999 -688 -1983 688
rect -2049 -700 -1983 -688
rect -1953 688 -1887 700
rect -1953 -688 -1937 688
rect -1903 -688 -1887 688
rect -1953 -700 -1887 -688
rect -1857 688 -1791 700
rect -1857 -688 -1841 688
rect -1807 -688 -1791 688
rect -1857 -700 -1791 -688
rect -1761 688 -1695 700
rect -1761 -688 -1745 688
rect -1711 -688 -1695 688
rect -1761 -700 -1695 -688
rect -1665 688 -1599 700
rect -1665 -688 -1649 688
rect -1615 -688 -1599 688
rect -1665 -700 -1599 -688
rect -1569 688 -1503 700
rect -1569 -688 -1553 688
rect -1519 -688 -1503 688
rect -1569 -700 -1503 -688
rect -1473 688 -1407 700
rect -1473 -688 -1457 688
rect -1423 -688 -1407 688
rect -1473 -700 -1407 -688
rect -1377 688 -1311 700
rect -1377 -688 -1361 688
rect -1327 -688 -1311 688
rect -1377 -700 -1311 -688
rect -1281 688 -1215 700
rect -1281 -688 -1265 688
rect -1231 -688 -1215 688
rect -1281 -700 -1215 -688
rect -1185 688 -1119 700
rect -1185 -688 -1169 688
rect -1135 -688 -1119 688
rect -1185 -700 -1119 -688
rect -1089 688 -1023 700
rect -1089 -688 -1073 688
rect -1039 -688 -1023 688
rect -1089 -700 -1023 -688
rect -993 688 -927 700
rect -993 -688 -977 688
rect -943 -688 -927 688
rect -993 -700 -927 -688
rect -897 688 -831 700
rect -897 -688 -881 688
rect -847 -688 -831 688
rect -897 -700 -831 -688
rect -801 688 -735 700
rect -801 -688 -785 688
rect -751 -688 -735 688
rect -801 -700 -735 -688
rect -705 688 -639 700
rect -705 -688 -689 688
rect -655 -688 -639 688
rect -705 -700 -639 -688
rect -609 688 -543 700
rect -609 -688 -593 688
rect -559 -688 -543 688
rect -609 -700 -543 -688
rect -513 688 -447 700
rect -513 -688 -497 688
rect -463 -688 -447 688
rect -513 -700 -447 -688
rect -417 688 -351 700
rect -417 -688 -401 688
rect -367 -688 -351 688
rect -417 -700 -351 -688
rect -321 688 -255 700
rect -321 -688 -305 688
rect -271 -688 -255 688
rect -321 -700 -255 -688
rect -225 688 -159 700
rect -225 -688 -209 688
rect -175 -688 -159 688
rect -225 -700 -159 -688
rect -129 688 -63 700
rect -129 -688 -113 688
rect -79 -688 -63 688
rect -129 -700 -63 -688
rect -33 688 33 700
rect -33 -688 -17 688
rect 17 -688 33 688
rect -33 -700 33 -688
rect 63 688 129 700
rect 63 -688 79 688
rect 113 -688 129 688
rect 63 -700 129 -688
rect 159 688 225 700
rect 159 -688 175 688
rect 209 -688 225 688
rect 159 -700 225 -688
rect 255 688 321 700
rect 255 -688 271 688
rect 305 -688 321 688
rect 255 -700 321 -688
rect 351 688 417 700
rect 351 -688 367 688
rect 401 -688 417 688
rect 351 -700 417 -688
rect 447 688 513 700
rect 447 -688 463 688
rect 497 -688 513 688
rect 447 -700 513 -688
rect 543 688 609 700
rect 543 -688 559 688
rect 593 -688 609 688
rect 543 -700 609 -688
rect 639 688 705 700
rect 639 -688 655 688
rect 689 -688 705 688
rect 639 -700 705 -688
rect 735 688 801 700
rect 735 -688 751 688
rect 785 -688 801 688
rect 735 -700 801 -688
rect 831 688 897 700
rect 831 -688 847 688
rect 881 -688 897 688
rect 831 -700 897 -688
rect 927 688 993 700
rect 927 -688 943 688
rect 977 -688 993 688
rect 927 -700 993 -688
rect 1023 688 1089 700
rect 1023 -688 1039 688
rect 1073 -688 1089 688
rect 1023 -700 1089 -688
rect 1119 688 1185 700
rect 1119 -688 1135 688
rect 1169 -688 1185 688
rect 1119 -700 1185 -688
rect 1215 688 1281 700
rect 1215 -688 1231 688
rect 1265 -688 1281 688
rect 1215 -700 1281 -688
rect 1311 688 1377 700
rect 1311 -688 1327 688
rect 1361 -688 1377 688
rect 1311 -700 1377 -688
rect 1407 688 1473 700
rect 1407 -688 1423 688
rect 1457 -688 1473 688
rect 1407 -700 1473 -688
rect 1503 688 1569 700
rect 1503 -688 1519 688
rect 1553 -688 1569 688
rect 1503 -700 1569 -688
rect 1599 688 1665 700
rect 1599 -688 1615 688
rect 1649 -688 1665 688
rect 1599 -700 1665 -688
rect 1695 688 1761 700
rect 1695 -688 1711 688
rect 1745 -688 1761 688
rect 1695 -700 1761 -688
rect 1791 688 1857 700
rect 1791 -688 1807 688
rect 1841 -688 1857 688
rect 1791 -700 1857 -688
rect 1887 688 1953 700
rect 1887 -688 1903 688
rect 1937 -688 1953 688
rect 1887 -700 1953 -688
rect 1983 688 2049 700
rect 1983 -688 1999 688
rect 2033 -688 2049 688
rect 1983 -700 2049 -688
rect 2079 688 2145 700
rect 2079 -688 2095 688
rect 2129 -688 2145 688
rect 2079 -700 2145 -688
rect 2175 688 2241 700
rect 2175 -688 2191 688
rect 2225 -688 2241 688
rect 2175 -700 2241 -688
rect 2271 688 2337 700
rect 2271 -688 2287 688
rect 2321 -688 2337 688
rect 2271 -700 2337 -688
rect 2367 688 2433 700
rect 2367 -688 2383 688
rect 2417 -688 2433 688
rect 2367 -700 2433 -688
rect 2463 688 2529 700
rect 2463 -688 2479 688
rect 2513 -688 2529 688
rect 2463 -700 2529 -688
rect 2559 688 2625 700
rect 2559 -688 2575 688
rect 2609 -688 2625 688
rect 2559 -700 2625 -688
rect 2655 688 2721 700
rect 2655 -688 2671 688
rect 2705 -688 2721 688
rect 2655 -700 2721 -688
rect 2751 688 2817 700
rect 2751 -688 2767 688
rect 2801 -688 2817 688
rect 2751 -700 2817 -688
rect 2847 688 2913 700
rect 2847 -688 2863 688
rect 2897 -688 2913 688
rect 2847 -700 2913 -688
rect 2943 688 3009 700
rect 2943 -688 2959 688
rect 2993 -688 3009 688
rect 2943 -700 3009 -688
rect 3039 688 3105 700
rect 3039 -688 3055 688
rect 3089 -688 3105 688
rect 3039 -700 3105 -688
rect 3135 688 3201 700
rect 3135 -688 3151 688
rect 3185 -688 3201 688
rect 3135 -700 3201 -688
rect 3231 688 3297 700
rect 3231 -688 3247 688
rect 3281 -688 3297 688
rect 3231 -700 3297 -688
rect 3327 688 3393 700
rect 3327 -688 3343 688
rect 3377 -688 3393 688
rect 3327 -700 3393 -688
rect 3423 688 3489 700
rect 3423 -688 3439 688
rect 3473 -688 3489 688
rect 3423 -700 3489 -688
rect 3519 688 3585 700
rect 3519 -688 3535 688
rect 3569 -688 3585 688
rect 3519 -700 3585 -688
rect 3615 688 3681 700
rect 3615 -688 3631 688
rect 3665 -688 3681 688
rect 3615 -700 3681 -688
rect 3711 688 3777 700
rect 3711 -688 3727 688
rect 3761 -688 3777 688
rect 3711 -700 3777 -688
rect 3807 688 3873 700
rect 3807 -688 3823 688
rect 3857 -688 3873 688
rect 3807 -700 3873 -688
rect 3903 688 3969 700
rect 3903 -688 3919 688
rect 3953 -688 3969 688
rect 3903 -700 3969 -688
rect 3999 688 4065 700
rect 3999 -688 4015 688
rect 4049 -688 4065 688
rect 3999 -700 4065 -688
rect 4095 688 4161 700
rect 4095 -688 4111 688
rect 4145 -688 4161 688
rect 4095 -700 4161 -688
rect 4191 688 4257 700
rect 4191 -688 4207 688
rect 4241 -688 4257 688
rect 4191 -700 4257 -688
rect 4287 688 4353 700
rect 4287 -688 4303 688
rect 4337 -688 4353 688
rect 4287 -700 4353 -688
rect 4383 688 4449 700
rect 4383 -688 4399 688
rect 4433 -688 4449 688
rect 4383 -700 4449 -688
rect 4479 688 4545 700
rect 4479 -688 4495 688
rect 4529 -688 4545 688
rect 4479 -700 4545 -688
rect 4575 688 4641 700
rect 4575 -688 4591 688
rect 4625 -688 4641 688
rect 4575 -700 4641 -688
rect 4671 688 4737 700
rect 4671 -688 4687 688
rect 4721 -688 4737 688
rect 4671 -700 4737 -688
rect 4767 688 4833 700
rect 4767 -688 4783 688
rect 4817 -688 4833 688
rect 4767 -700 4833 -688
rect 4863 688 4929 700
rect 4863 -688 4879 688
rect 4913 -688 4929 688
rect 4863 -700 4929 -688
rect 4959 688 5025 700
rect 4959 -688 4975 688
rect 5009 -688 5025 688
rect 4959 -700 5025 -688
rect 5055 688 5121 700
rect 5055 -688 5071 688
rect 5105 -688 5121 688
rect 5055 -700 5121 -688
rect 5151 688 5217 700
rect 5151 -688 5167 688
rect 5201 -688 5217 688
rect 5151 -700 5217 -688
rect 5247 688 5313 700
rect 5247 -688 5263 688
rect 5297 -688 5313 688
rect 5247 -700 5313 -688
rect 5343 688 5409 700
rect 5343 -688 5359 688
rect 5393 -688 5409 688
rect 5343 -700 5409 -688
rect 5439 688 5505 700
rect 5439 -688 5455 688
rect 5489 -688 5505 688
rect 5439 -700 5505 -688
rect 5535 688 5601 700
rect 5535 -688 5551 688
rect 5585 -688 5601 688
rect 5535 -700 5601 -688
rect 5631 688 5697 700
rect 5631 -688 5647 688
rect 5681 -688 5697 688
rect 5631 -700 5697 -688
rect 5727 688 5793 700
rect 5727 -688 5743 688
rect 5777 -688 5793 688
rect 5727 -700 5793 -688
rect 5823 688 5889 700
rect 5823 -688 5839 688
rect 5873 -688 5889 688
rect 5823 -700 5889 -688
rect 5919 688 5985 700
rect 5919 -688 5935 688
rect 5969 -688 5985 688
rect 5919 -700 5985 -688
rect 6015 688 6081 700
rect 6015 -688 6031 688
rect 6065 -688 6081 688
rect 6015 -700 6081 -688
rect 6111 688 6177 700
rect 6111 -688 6127 688
rect 6161 -688 6177 688
rect 6111 -700 6177 -688
rect 6207 688 6273 700
rect 6207 -688 6223 688
rect 6257 -688 6273 688
rect 6207 -700 6273 -688
rect 6303 688 6369 700
rect 6303 -688 6319 688
rect 6353 -688 6369 688
rect 6303 -700 6369 -688
rect 6399 688 6465 700
rect 6399 -688 6415 688
rect 6449 -688 6465 688
rect 6399 -700 6465 -688
rect 6495 688 6561 700
rect 6495 -688 6511 688
rect 6545 -688 6561 688
rect 6495 -700 6561 -688
rect 6591 688 6657 700
rect 6591 -688 6607 688
rect 6641 -688 6657 688
rect 6591 -700 6657 -688
rect 6687 688 6753 700
rect 6687 -688 6703 688
rect 6737 -688 6753 688
rect 6687 -700 6753 -688
rect 6783 688 6849 700
rect 6783 -688 6799 688
rect 6833 -688 6849 688
rect 6783 -700 6849 -688
rect 6879 688 6945 700
rect 6879 -688 6895 688
rect 6929 -688 6945 688
rect 6879 -700 6945 -688
rect 6975 688 7041 700
rect 6975 -688 6991 688
rect 7025 -688 7041 688
rect 6975 -700 7041 -688
rect 7071 688 7137 700
rect 7071 -688 7087 688
rect 7121 -688 7137 688
rect 7071 -700 7137 -688
rect 7167 688 7233 700
rect 7167 -688 7183 688
rect 7217 -688 7233 688
rect 7167 -700 7233 -688
rect 7263 688 7329 700
rect 7263 -688 7279 688
rect 7313 -688 7329 688
rect 7263 -700 7329 -688
rect 7359 688 7425 700
rect 7359 -688 7375 688
rect 7409 -688 7425 688
rect 7359 -700 7425 -688
rect 7455 688 7521 700
rect 7455 -688 7471 688
rect 7505 -688 7521 688
rect 7455 -700 7521 -688
rect 7551 688 7617 700
rect 7551 -688 7567 688
rect 7601 -688 7617 688
rect 7551 -700 7617 -688
rect 7647 688 7713 700
rect 7647 -688 7663 688
rect 7697 -688 7713 688
rect 7647 -700 7713 -688
rect 7743 688 7809 700
rect 7743 -688 7759 688
rect 7793 -688 7809 688
rect 7743 -700 7809 -688
rect 7839 688 7905 700
rect 7839 -688 7855 688
rect 7889 -688 7905 688
rect 7839 -700 7905 -688
rect 7935 688 8001 700
rect 7935 -688 7951 688
rect 7985 -688 8001 688
rect 7935 -700 8001 -688
rect 8031 688 8097 700
rect 8031 -688 8047 688
rect 8081 -688 8097 688
rect 8031 -700 8097 -688
rect 8127 688 8193 700
rect 8127 -688 8143 688
rect 8177 -688 8193 688
rect 8127 -700 8193 -688
rect 8223 688 8289 700
rect 8223 -688 8239 688
rect 8273 -688 8289 688
rect 8223 -700 8289 -688
rect 8319 688 8385 700
rect 8319 -688 8335 688
rect 8369 -688 8385 688
rect 8319 -700 8385 -688
rect 8415 688 8481 700
rect 8415 -688 8431 688
rect 8465 -688 8481 688
rect 8415 -700 8481 -688
rect 8511 688 8577 700
rect 8511 -688 8527 688
rect 8561 -688 8577 688
rect 8511 -700 8577 -688
rect 8607 688 8673 700
rect 8607 -688 8623 688
rect 8657 -688 8673 688
rect 8607 -700 8673 -688
rect 8703 688 8769 700
rect 8703 -688 8719 688
rect 8753 -688 8769 688
rect 8703 -700 8769 -688
rect 8799 688 8865 700
rect 8799 -688 8815 688
rect 8849 -688 8865 688
rect 8799 -700 8865 -688
rect 8895 688 8961 700
rect 8895 -688 8911 688
rect 8945 -688 8961 688
rect 8895 -700 8961 -688
rect 8991 688 9057 700
rect 8991 -688 9007 688
rect 9041 -688 9057 688
rect 8991 -700 9057 -688
rect 9087 688 9153 700
rect 9087 -688 9103 688
rect 9137 -688 9153 688
rect 9087 -700 9153 -688
rect 9183 688 9249 700
rect 9183 -688 9199 688
rect 9233 -688 9249 688
rect 9183 -700 9249 -688
rect 9279 688 9345 700
rect 9279 -688 9295 688
rect 9329 -688 9345 688
rect 9279 -700 9345 -688
rect 9375 688 9441 700
rect 9375 -688 9391 688
rect 9425 -688 9441 688
rect 9375 -700 9441 -688
rect 9471 688 9537 700
rect 9471 -688 9487 688
rect 9521 -688 9537 688
rect 9471 -700 9537 -688
rect 9567 688 9633 700
rect 9567 -688 9583 688
rect 9617 -688 9633 688
rect 9567 -700 9633 -688
rect 9663 688 9729 700
rect 9663 -688 9679 688
rect 9713 -688 9729 688
rect 9663 -700 9729 -688
rect 9759 688 9825 700
rect 9759 -688 9775 688
rect 9809 -688 9825 688
rect 9759 -700 9825 -688
rect 9855 688 9921 700
rect 9855 -688 9871 688
rect 9905 -688 9921 688
rect 9855 -700 9921 -688
rect 9951 688 10017 700
rect 9951 -688 9967 688
rect 10001 -688 10017 688
rect 9951 -700 10017 -688
rect 10047 688 10113 700
rect 10047 -688 10063 688
rect 10097 -688 10113 688
rect 10047 -700 10113 -688
rect 10143 688 10209 700
rect 10143 -688 10159 688
rect 10193 -688 10209 688
rect 10143 -700 10209 -688
rect 10239 688 10305 700
rect 10239 -688 10255 688
rect 10289 -688 10305 688
rect 10239 -700 10305 -688
rect 10335 688 10401 700
rect 10335 -688 10351 688
rect 10385 -688 10401 688
rect 10335 -700 10401 -688
rect 10431 688 10497 700
rect 10431 -688 10447 688
rect 10481 -688 10497 688
rect 10431 -700 10497 -688
rect 10527 688 10589 700
rect 10527 -688 10543 688
rect 10577 -688 10589 688
rect 10527 -700 10589 -688
<< pdiffc >>
rect -10577 -688 -10543 688
rect -10481 -688 -10447 688
rect -10385 -688 -10351 688
rect -10289 -688 -10255 688
rect -10193 -688 -10159 688
rect -10097 -688 -10063 688
rect -10001 -688 -9967 688
rect -9905 -688 -9871 688
rect -9809 -688 -9775 688
rect -9713 -688 -9679 688
rect -9617 -688 -9583 688
rect -9521 -688 -9487 688
rect -9425 -688 -9391 688
rect -9329 -688 -9295 688
rect -9233 -688 -9199 688
rect -9137 -688 -9103 688
rect -9041 -688 -9007 688
rect -8945 -688 -8911 688
rect -8849 -688 -8815 688
rect -8753 -688 -8719 688
rect -8657 -688 -8623 688
rect -8561 -688 -8527 688
rect -8465 -688 -8431 688
rect -8369 -688 -8335 688
rect -8273 -688 -8239 688
rect -8177 -688 -8143 688
rect -8081 -688 -8047 688
rect -7985 -688 -7951 688
rect -7889 -688 -7855 688
rect -7793 -688 -7759 688
rect -7697 -688 -7663 688
rect -7601 -688 -7567 688
rect -7505 -688 -7471 688
rect -7409 -688 -7375 688
rect -7313 -688 -7279 688
rect -7217 -688 -7183 688
rect -7121 -688 -7087 688
rect -7025 -688 -6991 688
rect -6929 -688 -6895 688
rect -6833 -688 -6799 688
rect -6737 -688 -6703 688
rect -6641 -688 -6607 688
rect -6545 -688 -6511 688
rect -6449 -688 -6415 688
rect -6353 -688 -6319 688
rect -6257 -688 -6223 688
rect -6161 -688 -6127 688
rect -6065 -688 -6031 688
rect -5969 -688 -5935 688
rect -5873 -688 -5839 688
rect -5777 -688 -5743 688
rect -5681 -688 -5647 688
rect -5585 -688 -5551 688
rect -5489 -688 -5455 688
rect -5393 -688 -5359 688
rect -5297 -688 -5263 688
rect -5201 -688 -5167 688
rect -5105 -688 -5071 688
rect -5009 -688 -4975 688
rect -4913 -688 -4879 688
rect -4817 -688 -4783 688
rect -4721 -688 -4687 688
rect -4625 -688 -4591 688
rect -4529 -688 -4495 688
rect -4433 -688 -4399 688
rect -4337 -688 -4303 688
rect -4241 -688 -4207 688
rect -4145 -688 -4111 688
rect -4049 -688 -4015 688
rect -3953 -688 -3919 688
rect -3857 -688 -3823 688
rect -3761 -688 -3727 688
rect -3665 -688 -3631 688
rect -3569 -688 -3535 688
rect -3473 -688 -3439 688
rect -3377 -688 -3343 688
rect -3281 -688 -3247 688
rect -3185 -688 -3151 688
rect -3089 -688 -3055 688
rect -2993 -688 -2959 688
rect -2897 -688 -2863 688
rect -2801 -688 -2767 688
rect -2705 -688 -2671 688
rect -2609 -688 -2575 688
rect -2513 -688 -2479 688
rect -2417 -688 -2383 688
rect -2321 -688 -2287 688
rect -2225 -688 -2191 688
rect -2129 -688 -2095 688
rect -2033 -688 -1999 688
rect -1937 -688 -1903 688
rect -1841 -688 -1807 688
rect -1745 -688 -1711 688
rect -1649 -688 -1615 688
rect -1553 -688 -1519 688
rect -1457 -688 -1423 688
rect -1361 -688 -1327 688
rect -1265 -688 -1231 688
rect -1169 -688 -1135 688
rect -1073 -688 -1039 688
rect -977 -688 -943 688
rect -881 -688 -847 688
rect -785 -688 -751 688
rect -689 -688 -655 688
rect -593 -688 -559 688
rect -497 -688 -463 688
rect -401 -688 -367 688
rect -305 -688 -271 688
rect -209 -688 -175 688
rect -113 -688 -79 688
rect -17 -688 17 688
rect 79 -688 113 688
rect 175 -688 209 688
rect 271 -688 305 688
rect 367 -688 401 688
rect 463 -688 497 688
rect 559 -688 593 688
rect 655 -688 689 688
rect 751 -688 785 688
rect 847 -688 881 688
rect 943 -688 977 688
rect 1039 -688 1073 688
rect 1135 -688 1169 688
rect 1231 -688 1265 688
rect 1327 -688 1361 688
rect 1423 -688 1457 688
rect 1519 -688 1553 688
rect 1615 -688 1649 688
rect 1711 -688 1745 688
rect 1807 -688 1841 688
rect 1903 -688 1937 688
rect 1999 -688 2033 688
rect 2095 -688 2129 688
rect 2191 -688 2225 688
rect 2287 -688 2321 688
rect 2383 -688 2417 688
rect 2479 -688 2513 688
rect 2575 -688 2609 688
rect 2671 -688 2705 688
rect 2767 -688 2801 688
rect 2863 -688 2897 688
rect 2959 -688 2993 688
rect 3055 -688 3089 688
rect 3151 -688 3185 688
rect 3247 -688 3281 688
rect 3343 -688 3377 688
rect 3439 -688 3473 688
rect 3535 -688 3569 688
rect 3631 -688 3665 688
rect 3727 -688 3761 688
rect 3823 -688 3857 688
rect 3919 -688 3953 688
rect 4015 -688 4049 688
rect 4111 -688 4145 688
rect 4207 -688 4241 688
rect 4303 -688 4337 688
rect 4399 -688 4433 688
rect 4495 -688 4529 688
rect 4591 -688 4625 688
rect 4687 -688 4721 688
rect 4783 -688 4817 688
rect 4879 -688 4913 688
rect 4975 -688 5009 688
rect 5071 -688 5105 688
rect 5167 -688 5201 688
rect 5263 -688 5297 688
rect 5359 -688 5393 688
rect 5455 -688 5489 688
rect 5551 -688 5585 688
rect 5647 -688 5681 688
rect 5743 -688 5777 688
rect 5839 -688 5873 688
rect 5935 -688 5969 688
rect 6031 -688 6065 688
rect 6127 -688 6161 688
rect 6223 -688 6257 688
rect 6319 -688 6353 688
rect 6415 -688 6449 688
rect 6511 -688 6545 688
rect 6607 -688 6641 688
rect 6703 -688 6737 688
rect 6799 -688 6833 688
rect 6895 -688 6929 688
rect 6991 -688 7025 688
rect 7087 -688 7121 688
rect 7183 -688 7217 688
rect 7279 -688 7313 688
rect 7375 -688 7409 688
rect 7471 -688 7505 688
rect 7567 -688 7601 688
rect 7663 -688 7697 688
rect 7759 -688 7793 688
rect 7855 -688 7889 688
rect 7951 -688 7985 688
rect 8047 -688 8081 688
rect 8143 -688 8177 688
rect 8239 -688 8273 688
rect 8335 -688 8369 688
rect 8431 -688 8465 688
rect 8527 -688 8561 688
rect 8623 -688 8657 688
rect 8719 -688 8753 688
rect 8815 -688 8849 688
rect 8911 -688 8945 688
rect 9007 -688 9041 688
rect 9103 -688 9137 688
rect 9199 -688 9233 688
rect 9295 -688 9329 688
rect 9391 -688 9425 688
rect 9487 -688 9521 688
rect 9583 -688 9617 688
rect 9679 -688 9713 688
rect 9775 -688 9809 688
rect 9871 -688 9905 688
rect 9967 -688 10001 688
rect 10063 -688 10097 688
rect 10159 -688 10193 688
rect 10255 -688 10289 688
rect 10351 -688 10385 688
rect 10447 -688 10481 688
rect 10543 -688 10577 688
<< nsubdiff >>
rect -10691 849 -10595 883
rect 10595 849 10691 883
rect -10691 787 -10657 849
rect 10657 787 10691 849
rect -10691 -849 -10657 -787
rect 10657 -849 10691 -787
rect -10691 -883 -10595 -849
rect 10595 -883 10691 -849
<< nsubdiffcont >>
rect -10595 849 10595 883
rect -10691 -787 -10657 787
rect 10657 -787 10691 787
rect -10595 -883 10595 -849
<< poly >>
rect -10449 781 -10383 797
rect -10449 747 -10433 781
rect -10399 747 -10383 781
rect -10449 731 -10383 747
rect -10257 781 -10191 797
rect -10257 747 -10241 781
rect -10207 747 -10191 781
rect -10257 731 -10191 747
rect -10065 781 -9999 797
rect -10065 747 -10049 781
rect -10015 747 -9999 781
rect -10065 731 -9999 747
rect -9873 781 -9807 797
rect -9873 747 -9857 781
rect -9823 747 -9807 781
rect -9873 731 -9807 747
rect -9681 781 -9615 797
rect -9681 747 -9665 781
rect -9631 747 -9615 781
rect -9681 731 -9615 747
rect -9489 781 -9423 797
rect -9489 747 -9473 781
rect -9439 747 -9423 781
rect -9489 731 -9423 747
rect -9297 781 -9231 797
rect -9297 747 -9281 781
rect -9247 747 -9231 781
rect -9297 731 -9231 747
rect -9105 781 -9039 797
rect -9105 747 -9089 781
rect -9055 747 -9039 781
rect -9105 731 -9039 747
rect -8913 781 -8847 797
rect -8913 747 -8897 781
rect -8863 747 -8847 781
rect -8913 731 -8847 747
rect -8721 781 -8655 797
rect -8721 747 -8705 781
rect -8671 747 -8655 781
rect -8721 731 -8655 747
rect -8529 781 -8463 797
rect -8529 747 -8513 781
rect -8479 747 -8463 781
rect -8529 731 -8463 747
rect -8337 781 -8271 797
rect -8337 747 -8321 781
rect -8287 747 -8271 781
rect -8337 731 -8271 747
rect -8145 781 -8079 797
rect -8145 747 -8129 781
rect -8095 747 -8079 781
rect -8145 731 -8079 747
rect -7953 781 -7887 797
rect -7953 747 -7937 781
rect -7903 747 -7887 781
rect -7953 731 -7887 747
rect -7761 781 -7695 797
rect -7761 747 -7745 781
rect -7711 747 -7695 781
rect -7761 731 -7695 747
rect -7569 781 -7503 797
rect -7569 747 -7553 781
rect -7519 747 -7503 781
rect -7569 731 -7503 747
rect -7377 781 -7311 797
rect -7377 747 -7361 781
rect -7327 747 -7311 781
rect -7377 731 -7311 747
rect -7185 781 -7119 797
rect -7185 747 -7169 781
rect -7135 747 -7119 781
rect -7185 731 -7119 747
rect -6993 781 -6927 797
rect -6993 747 -6977 781
rect -6943 747 -6927 781
rect -6993 731 -6927 747
rect -6801 781 -6735 797
rect -6801 747 -6785 781
rect -6751 747 -6735 781
rect -6801 731 -6735 747
rect -6609 781 -6543 797
rect -6609 747 -6593 781
rect -6559 747 -6543 781
rect -6609 731 -6543 747
rect -6417 781 -6351 797
rect -6417 747 -6401 781
rect -6367 747 -6351 781
rect -6417 731 -6351 747
rect -6225 781 -6159 797
rect -6225 747 -6209 781
rect -6175 747 -6159 781
rect -6225 731 -6159 747
rect -6033 781 -5967 797
rect -6033 747 -6017 781
rect -5983 747 -5967 781
rect -6033 731 -5967 747
rect -5841 781 -5775 797
rect -5841 747 -5825 781
rect -5791 747 -5775 781
rect -5841 731 -5775 747
rect -5649 781 -5583 797
rect -5649 747 -5633 781
rect -5599 747 -5583 781
rect -5649 731 -5583 747
rect -5457 781 -5391 797
rect -5457 747 -5441 781
rect -5407 747 -5391 781
rect -5457 731 -5391 747
rect -5265 781 -5199 797
rect -5265 747 -5249 781
rect -5215 747 -5199 781
rect -5265 731 -5199 747
rect -5073 781 -5007 797
rect -5073 747 -5057 781
rect -5023 747 -5007 781
rect -5073 731 -5007 747
rect -4881 781 -4815 797
rect -4881 747 -4865 781
rect -4831 747 -4815 781
rect -4881 731 -4815 747
rect -4689 781 -4623 797
rect -4689 747 -4673 781
rect -4639 747 -4623 781
rect -4689 731 -4623 747
rect -4497 781 -4431 797
rect -4497 747 -4481 781
rect -4447 747 -4431 781
rect -4497 731 -4431 747
rect -4305 781 -4239 797
rect -4305 747 -4289 781
rect -4255 747 -4239 781
rect -4305 731 -4239 747
rect -4113 781 -4047 797
rect -4113 747 -4097 781
rect -4063 747 -4047 781
rect -4113 731 -4047 747
rect -3921 781 -3855 797
rect -3921 747 -3905 781
rect -3871 747 -3855 781
rect -3921 731 -3855 747
rect -3729 781 -3663 797
rect -3729 747 -3713 781
rect -3679 747 -3663 781
rect -3729 731 -3663 747
rect -3537 781 -3471 797
rect -3537 747 -3521 781
rect -3487 747 -3471 781
rect -3537 731 -3471 747
rect -3345 781 -3279 797
rect -3345 747 -3329 781
rect -3295 747 -3279 781
rect -3345 731 -3279 747
rect -3153 781 -3087 797
rect -3153 747 -3137 781
rect -3103 747 -3087 781
rect -3153 731 -3087 747
rect -2961 781 -2895 797
rect -2961 747 -2945 781
rect -2911 747 -2895 781
rect -2961 731 -2895 747
rect -2769 781 -2703 797
rect -2769 747 -2753 781
rect -2719 747 -2703 781
rect -2769 731 -2703 747
rect -2577 781 -2511 797
rect -2577 747 -2561 781
rect -2527 747 -2511 781
rect -2577 731 -2511 747
rect -2385 781 -2319 797
rect -2385 747 -2369 781
rect -2335 747 -2319 781
rect -2385 731 -2319 747
rect -2193 781 -2127 797
rect -2193 747 -2177 781
rect -2143 747 -2127 781
rect -2193 731 -2127 747
rect -2001 781 -1935 797
rect -2001 747 -1985 781
rect -1951 747 -1935 781
rect -2001 731 -1935 747
rect -1809 781 -1743 797
rect -1809 747 -1793 781
rect -1759 747 -1743 781
rect -1809 731 -1743 747
rect -1617 781 -1551 797
rect -1617 747 -1601 781
rect -1567 747 -1551 781
rect -1617 731 -1551 747
rect -1425 781 -1359 797
rect -1425 747 -1409 781
rect -1375 747 -1359 781
rect -1425 731 -1359 747
rect -1233 781 -1167 797
rect -1233 747 -1217 781
rect -1183 747 -1167 781
rect -1233 731 -1167 747
rect -1041 781 -975 797
rect -1041 747 -1025 781
rect -991 747 -975 781
rect -1041 731 -975 747
rect -849 781 -783 797
rect -849 747 -833 781
rect -799 747 -783 781
rect -849 731 -783 747
rect -657 781 -591 797
rect -657 747 -641 781
rect -607 747 -591 781
rect -657 731 -591 747
rect -465 781 -399 797
rect -465 747 -449 781
rect -415 747 -399 781
rect -465 731 -399 747
rect -273 781 -207 797
rect -273 747 -257 781
rect -223 747 -207 781
rect -273 731 -207 747
rect -81 781 -15 797
rect -81 747 -65 781
rect -31 747 -15 781
rect -81 731 -15 747
rect 111 781 177 797
rect 111 747 127 781
rect 161 747 177 781
rect 111 731 177 747
rect 303 781 369 797
rect 303 747 319 781
rect 353 747 369 781
rect 303 731 369 747
rect 495 781 561 797
rect 495 747 511 781
rect 545 747 561 781
rect 495 731 561 747
rect 687 781 753 797
rect 687 747 703 781
rect 737 747 753 781
rect 687 731 753 747
rect 879 781 945 797
rect 879 747 895 781
rect 929 747 945 781
rect 879 731 945 747
rect 1071 781 1137 797
rect 1071 747 1087 781
rect 1121 747 1137 781
rect 1071 731 1137 747
rect 1263 781 1329 797
rect 1263 747 1279 781
rect 1313 747 1329 781
rect 1263 731 1329 747
rect 1455 781 1521 797
rect 1455 747 1471 781
rect 1505 747 1521 781
rect 1455 731 1521 747
rect 1647 781 1713 797
rect 1647 747 1663 781
rect 1697 747 1713 781
rect 1647 731 1713 747
rect 1839 781 1905 797
rect 1839 747 1855 781
rect 1889 747 1905 781
rect 1839 731 1905 747
rect 2031 781 2097 797
rect 2031 747 2047 781
rect 2081 747 2097 781
rect 2031 731 2097 747
rect 2223 781 2289 797
rect 2223 747 2239 781
rect 2273 747 2289 781
rect 2223 731 2289 747
rect 2415 781 2481 797
rect 2415 747 2431 781
rect 2465 747 2481 781
rect 2415 731 2481 747
rect 2607 781 2673 797
rect 2607 747 2623 781
rect 2657 747 2673 781
rect 2607 731 2673 747
rect 2799 781 2865 797
rect 2799 747 2815 781
rect 2849 747 2865 781
rect 2799 731 2865 747
rect 2991 781 3057 797
rect 2991 747 3007 781
rect 3041 747 3057 781
rect 2991 731 3057 747
rect 3183 781 3249 797
rect 3183 747 3199 781
rect 3233 747 3249 781
rect 3183 731 3249 747
rect 3375 781 3441 797
rect 3375 747 3391 781
rect 3425 747 3441 781
rect 3375 731 3441 747
rect 3567 781 3633 797
rect 3567 747 3583 781
rect 3617 747 3633 781
rect 3567 731 3633 747
rect 3759 781 3825 797
rect 3759 747 3775 781
rect 3809 747 3825 781
rect 3759 731 3825 747
rect 3951 781 4017 797
rect 3951 747 3967 781
rect 4001 747 4017 781
rect 3951 731 4017 747
rect 4143 781 4209 797
rect 4143 747 4159 781
rect 4193 747 4209 781
rect 4143 731 4209 747
rect 4335 781 4401 797
rect 4335 747 4351 781
rect 4385 747 4401 781
rect 4335 731 4401 747
rect 4527 781 4593 797
rect 4527 747 4543 781
rect 4577 747 4593 781
rect 4527 731 4593 747
rect 4719 781 4785 797
rect 4719 747 4735 781
rect 4769 747 4785 781
rect 4719 731 4785 747
rect 4911 781 4977 797
rect 4911 747 4927 781
rect 4961 747 4977 781
rect 4911 731 4977 747
rect 5103 781 5169 797
rect 5103 747 5119 781
rect 5153 747 5169 781
rect 5103 731 5169 747
rect 5295 781 5361 797
rect 5295 747 5311 781
rect 5345 747 5361 781
rect 5295 731 5361 747
rect 5487 781 5553 797
rect 5487 747 5503 781
rect 5537 747 5553 781
rect 5487 731 5553 747
rect 5679 781 5745 797
rect 5679 747 5695 781
rect 5729 747 5745 781
rect 5679 731 5745 747
rect 5871 781 5937 797
rect 5871 747 5887 781
rect 5921 747 5937 781
rect 5871 731 5937 747
rect 6063 781 6129 797
rect 6063 747 6079 781
rect 6113 747 6129 781
rect 6063 731 6129 747
rect 6255 781 6321 797
rect 6255 747 6271 781
rect 6305 747 6321 781
rect 6255 731 6321 747
rect 6447 781 6513 797
rect 6447 747 6463 781
rect 6497 747 6513 781
rect 6447 731 6513 747
rect 6639 781 6705 797
rect 6639 747 6655 781
rect 6689 747 6705 781
rect 6639 731 6705 747
rect 6831 781 6897 797
rect 6831 747 6847 781
rect 6881 747 6897 781
rect 6831 731 6897 747
rect 7023 781 7089 797
rect 7023 747 7039 781
rect 7073 747 7089 781
rect 7023 731 7089 747
rect 7215 781 7281 797
rect 7215 747 7231 781
rect 7265 747 7281 781
rect 7215 731 7281 747
rect 7407 781 7473 797
rect 7407 747 7423 781
rect 7457 747 7473 781
rect 7407 731 7473 747
rect 7599 781 7665 797
rect 7599 747 7615 781
rect 7649 747 7665 781
rect 7599 731 7665 747
rect 7791 781 7857 797
rect 7791 747 7807 781
rect 7841 747 7857 781
rect 7791 731 7857 747
rect 7983 781 8049 797
rect 7983 747 7999 781
rect 8033 747 8049 781
rect 7983 731 8049 747
rect 8175 781 8241 797
rect 8175 747 8191 781
rect 8225 747 8241 781
rect 8175 731 8241 747
rect 8367 781 8433 797
rect 8367 747 8383 781
rect 8417 747 8433 781
rect 8367 731 8433 747
rect 8559 781 8625 797
rect 8559 747 8575 781
rect 8609 747 8625 781
rect 8559 731 8625 747
rect 8751 781 8817 797
rect 8751 747 8767 781
rect 8801 747 8817 781
rect 8751 731 8817 747
rect 8943 781 9009 797
rect 8943 747 8959 781
rect 8993 747 9009 781
rect 8943 731 9009 747
rect 9135 781 9201 797
rect 9135 747 9151 781
rect 9185 747 9201 781
rect 9135 731 9201 747
rect 9327 781 9393 797
rect 9327 747 9343 781
rect 9377 747 9393 781
rect 9327 731 9393 747
rect 9519 781 9585 797
rect 9519 747 9535 781
rect 9569 747 9585 781
rect 9519 731 9585 747
rect 9711 781 9777 797
rect 9711 747 9727 781
rect 9761 747 9777 781
rect 9711 731 9777 747
rect 9903 781 9969 797
rect 9903 747 9919 781
rect 9953 747 9969 781
rect 9903 731 9969 747
rect 10095 781 10161 797
rect 10095 747 10111 781
rect 10145 747 10161 781
rect 10095 731 10161 747
rect 10287 781 10353 797
rect 10287 747 10303 781
rect 10337 747 10353 781
rect 10287 731 10353 747
rect 10479 781 10545 797
rect 10479 747 10495 781
rect 10529 747 10545 781
rect 10479 731 10545 747
rect -10527 700 -10497 726
rect -10431 700 -10401 731
rect -10335 700 -10305 726
rect -10239 700 -10209 731
rect -10143 700 -10113 726
rect -10047 700 -10017 731
rect -9951 700 -9921 726
rect -9855 700 -9825 731
rect -9759 700 -9729 726
rect -9663 700 -9633 731
rect -9567 700 -9537 726
rect -9471 700 -9441 731
rect -9375 700 -9345 726
rect -9279 700 -9249 731
rect -9183 700 -9153 726
rect -9087 700 -9057 731
rect -8991 700 -8961 726
rect -8895 700 -8865 731
rect -8799 700 -8769 726
rect -8703 700 -8673 731
rect -8607 700 -8577 726
rect -8511 700 -8481 731
rect -8415 700 -8385 726
rect -8319 700 -8289 731
rect -8223 700 -8193 726
rect -8127 700 -8097 731
rect -8031 700 -8001 726
rect -7935 700 -7905 731
rect -7839 700 -7809 726
rect -7743 700 -7713 731
rect -7647 700 -7617 726
rect -7551 700 -7521 731
rect -7455 700 -7425 726
rect -7359 700 -7329 731
rect -7263 700 -7233 726
rect -7167 700 -7137 731
rect -7071 700 -7041 726
rect -6975 700 -6945 731
rect -6879 700 -6849 726
rect -6783 700 -6753 731
rect -6687 700 -6657 726
rect -6591 700 -6561 731
rect -6495 700 -6465 726
rect -6399 700 -6369 731
rect -6303 700 -6273 726
rect -6207 700 -6177 731
rect -6111 700 -6081 726
rect -6015 700 -5985 731
rect -5919 700 -5889 726
rect -5823 700 -5793 731
rect -5727 700 -5697 726
rect -5631 700 -5601 731
rect -5535 700 -5505 726
rect -5439 700 -5409 731
rect -5343 700 -5313 726
rect -5247 700 -5217 731
rect -5151 700 -5121 726
rect -5055 700 -5025 731
rect -4959 700 -4929 726
rect -4863 700 -4833 731
rect -4767 700 -4737 726
rect -4671 700 -4641 731
rect -4575 700 -4545 726
rect -4479 700 -4449 731
rect -4383 700 -4353 726
rect -4287 700 -4257 731
rect -4191 700 -4161 726
rect -4095 700 -4065 731
rect -3999 700 -3969 726
rect -3903 700 -3873 731
rect -3807 700 -3777 726
rect -3711 700 -3681 731
rect -3615 700 -3585 726
rect -3519 700 -3489 731
rect -3423 700 -3393 726
rect -3327 700 -3297 731
rect -3231 700 -3201 726
rect -3135 700 -3105 731
rect -3039 700 -3009 726
rect -2943 700 -2913 731
rect -2847 700 -2817 726
rect -2751 700 -2721 731
rect -2655 700 -2625 726
rect -2559 700 -2529 731
rect -2463 700 -2433 726
rect -2367 700 -2337 731
rect -2271 700 -2241 726
rect -2175 700 -2145 731
rect -2079 700 -2049 726
rect -1983 700 -1953 731
rect -1887 700 -1857 726
rect -1791 700 -1761 731
rect -1695 700 -1665 726
rect -1599 700 -1569 731
rect -1503 700 -1473 726
rect -1407 700 -1377 731
rect -1311 700 -1281 726
rect -1215 700 -1185 731
rect -1119 700 -1089 726
rect -1023 700 -993 731
rect -927 700 -897 726
rect -831 700 -801 731
rect -735 700 -705 726
rect -639 700 -609 731
rect -543 700 -513 726
rect -447 700 -417 731
rect -351 700 -321 726
rect -255 700 -225 731
rect -159 700 -129 726
rect -63 700 -33 731
rect 33 700 63 726
rect 129 700 159 731
rect 225 700 255 726
rect 321 700 351 731
rect 417 700 447 726
rect 513 700 543 731
rect 609 700 639 726
rect 705 700 735 731
rect 801 700 831 726
rect 897 700 927 731
rect 993 700 1023 726
rect 1089 700 1119 731
rect 1185 700 1215 726
rect 1281 700 1311 731
rect 1377 700 1407 726
rect 1473 700 1503 731
rect 1569 700 1599 726
rect 1665 700 1695 731
rect 1761 700 1791 726
rect 1857 700 1887 731
rect 1953 700 1983 726
rect 2049 700 2079 731
rect 2145 700 2175 726
rect 2241 700 2271 731
rect 2337 700 2367 726
rect 2433 700 2463 731
rect 2529 700 2559 726
rect 2625 700 2655 731
rect 2721 700 2751 726
rect 2817 700 2847 731
rect 2913 700 2943 726
rect 3009 700 3039 731
rect 3105 700 3135 726
rect 3201 700 3231 731
rect 3297 700 3327 726
rect 3393 700 3423 731
rect 3489 700 3519 726
rect 3585 700 3615 731
rect 3681 700 3711 726
rect 3777 700 3807 731
rect 3873 700 3903 726
rect 3969 700 3999 731
rect 4065 700 4095 726
rect 4161 700 4191 731
rect 4257 700 4287 726
rect 4353 700 4383 731
rect 4449 700 4479 726
rect 4545 700 4575 731
rect 4641 700 4671 726
rect 4737 700 4767 731
rect 4833 700 4863 726
rect 4929 700 4959 731
rect 5025 700 5055 726
rect 5121 700 5151 731
rect 5217 700 5247 726
rect 5313 700 5343 731
rect 5409 700 5439 726
rect 5505 700 5535 731
rect 5601 700 5631 726
rect 5697 700 5727 731
rect 5793 700 5823 726
rect 5889 700 5919 731
rect 5985 700 6015 726
rect 6081 700 6111 731
rect 6177 700 6207 726
rect 6273 700 6303 731
rect 6369 700 6399 726
rect 6465 700 6495 731
rect 6561 700 6591 726
rect 6657 700 6687 731
rect 6753 700 6783 726
rect 6849 700 6879 731
rect 6945 700 6975 726
rect 7041 700 7071 731
rect 7137 700 7167 726
rect 7233 700 7263 731
rect 7329 700 7359 726
rect 7425 700 7455 731
rect 7521 700 7551 726
rect 7617 700 7647 731
rect 7713 700 7743 726
rect 7809 700 7839 731
rect 7905 700 7935 726
rect 8001 700 8031 731
rect 8097 700 8127 726
rect 8193 700 8223 731
rect 8289 700 8319 726
rect 8385 700 8415 731
rect 8481 700 8511 726
rect 8577 700 8607 731
rect 8673 700 8703 726
rect 8769 700 8799 731
rect 8865 700 8895 726
rect 8961 700 8991 731
rect 9057 700 9087 726
rect 9153 700 9183 731
rect 9249 700 9279 726
rect 9345 700 9375 731
rect 9441 700 9471 726
rect 9537 700 9567 731
rect 9633 700 9663 726
rect 9729 700 9759 731
rect 9825 700 9855 726
rect 9921 700 9951 731
rect 10017 700 10047 726
rect 10113 700 10143 731
rect 10209 700 10239 726
rect 10305 700 10335 731
rect 10401 700 10431 726
rect 10497 700 10527 731
rect -10527 -731 -10497 -700
rect -10431 -726 -10401 -700
rect -10335 -731 -10305 -700
rect -10239 -726 -10209 -700
rect -10143 -731 -10113 -700
rect -10047 -726 -10017 -700
rect -9951 -731 -9921 -700
rect -9855 -726 -9825 -700
rect -9759 -731 -9729 -700
rect -9663 -726 -9633 -700
rect -9567 -731 -9537 -700
rect -9471 -726 -9441 -700
rect -9375 -731 -9345 -700
rect -9279 -726 -9249 -700
rect -9183 -731 -9153 -700
rect -9087 -726 -9057 -700
rect -8991 -731 -8961 -700
rect -8895 -726 -8865 -700
rect -8799 -731 -8769 -700
rect -8703 -726 -8673 -700
rect -8607 -731 -8577 -700
rect -8511 -726 -8481 -700
rect -8415 -731 -8385 -700
rect -8319 -726 -8289 -700
rect -8223 -731 -8193 -700
rect -8127 -726 -8097 -700
rect -8031 -731 -8001 -700
rect -7935 -726 -7905 -700
rect -7839 -731 -7809 -700
rect -7743 -726 -7713 -700
rect -7647 -731 -7617 -700
rect -7551 -726 -7521 -700
rect -7455 -731 -7425 -700
rect -7359 -726 -7329 -700
rect -7263 -731 -7233 -700
rect -7167 -726 -7137 -700
rect -7071 -731 -7041 -700
rect -6975 -726 -6945 -700
rect -6879 -731 -6849 -700
rect -6783 -726 -6753 -700
rect -6687 -731 -6657 -700
rect -6591 -726 -6561 -700
rect -6495 -731 -6465 -700
rect -6399 -726 -6369 -700
rect -6303 -731 -6273 -700
rect -6207 -726 -6177 -700
rect -6111 -731 -6081 -700
rect -6015 -726 -5985 -700
rect -5919 -731 -5889 -700
rect -5823 -726 -5793 -700
rect -5727 -731 -5697 -700
rect -5631 -726 -5601 -700
rect -5535 -731 -5505 -700
rect -5439 -726 -5409 -700
rect -5343 -731 -5313 -700
rect -5247 -726 -5217 -700
rect -5151 -731 -5121 -700
rect -5055 -726 -5025 -700
rect -4959 -731 -4929 -700
rect -4863 -726 -4833 -700
rect -4767 -731 -4737 -700
rect -4671 -726 -4641 -700
rect -4575 -731 -4545 -700
rect -4479 -726 -4449 -700
rect -4383 -731 -4353 -700
rect -4287 -726 -4257 -700
rect -4191 -731 -4161 -700
rect -4095 -726 -4065 -700
rect -3999 -731 -3969 -700
rect -3903 -726 -3873 -700
rect -3807 -731 -3777 -700
rect -3711 -726 -3681 -700
rect -3615 -731 -3585 -700
rect -3519 -726 -3489 -700
rect -3423 -731 -3393 -700
rect -3327 -726 -3297 -700
rect -3231 -731 -3201 -700
rect -3135 -726 -3105 -700
rect -3039 -731 -3009 -700
rect -2943 -726 -2913 -700
rect -2847 -731 -2817 -700
rect -2751 -726 -2721 -700
rect -2655 -731 -2625 -700
rect -2559 -726 -2529 -700
rect -2463 -731 -2433 -700
rect -2367 -726 -2337 -700
rect -2271 -731 -2241 -700
rect -2175 -726 -2145 -700
rect -2079 -731 -2049 -700
rect -1983 -726 -1953 -700
rect -1887 -731 -1857 -700
rect -1791 -726 -1761 -700
rect -1695 -731 -1665 -700
rect -1599 -726 -1569 -700
rect -1503 -731 -1473 -700
rect -1407 -726 -1377 -700
rect -1311 -731 -1281 -700
rect -1215 -726 -1185 -700
rect -1119 -731 -1089 -700
rect -1023 -726 -993 -700
rect -927 -731 -897 -700
rect -831 -726 -801 -700
rect -735 -731 -705 -700
rect -639 -726 -609 -700
rect -543 -731 -513 -700
rect -447 -726 -417 -700
rect -351 -731 -321 -700
rect -255 -726 -225 -700
rect -159 -731 -129 -700
rect -63 -726 -33 -700
rect 33 -731 63 -700
rect 129 -726 159 -700
rect 225 -731 255 -700
rect 321 -726 351 -700
rect 417 -731 447 -700
rect 513 -726 543 -700
rect 609 -731 639 -700
rect 705 -726 735 -700
rect 801 -731 831 -700
rect 897 -726 927 -700
rect 993 -731 1023 -700
rect 1089 -726 1119 -700
rect 1185 -731 1215 -700
rect 1281 -726 1311 -700
rect 1377 -731 1407 -700
rect 1473 -726 1503 -700
rect 1569 -731 1599 -700
rect 1665 -726 1695 -700
rect 1761 -731 1791 -700
rect 1857 -726 1887 -700
rect 1953 -731 1983 -700
rect 2049 -726 2079 -700
rect 2145 -731 2175 -700
rect 2241 -726 2271 -700
rect 2337 -731 2367 -700
rect 2433 -726 2463 -700
rect 2529 -731 2559 -700
rect 2625 -726 2655 -700
rect 2721 -731 2751 -700
rect 2817 -726 2847 -700
rect 2913 -731 2943 -700
rect 3009 -726 3039 -700
rect 3105 -731 3135 -700
rect 3201 -726 3231 -700
rect 3297 -731 3327 -700
rect 3393 -726 3423 -700
rect 3489 -731 3519 -700
rect 3585 -726 3615 -700
rect 3681 -731 3711 -700
rect 3777 -726 3807 -700
rect 3873 -731 3903 -700
rect 3969 -726 3999 -700
rect 4065 -731 4095 -700
rect 4161 -726 4191 -700
rect 4257 -731 4287 -700
rect 4353 -726 4383 -700
rect 4449 -731 4479 -700
rect 4545 -726 4575 -700
rect 4641 -731 4671 -700
rect 4737 -726 4767 -700
rect 4833 -731 4863 -700
rect 4929 -726 4959 -700
rect 5025 -731 5055 -700
rect 5121 -726 5151 -700
rect 5217 -731 5247 -700
rect 5313 -726 5343 -700
rect 5409 -731 5439 -700
rect 5505 -726 5535 -700
rect 5601 -731 5631 -700
rect 5697 -726 5727 -700
rect 5793 -731 5823 -700
rect 5889 -726 5919 -700
rect 5985 -731 6015 -700
rect 6081 -726 6111 -700
rect 6177 -731 6207 -700
rect 6273 -726 6303 -700
rect 6369 -731 6399 -700
rect 6465 -726 6495 -700
rect 6561 -731 6591 -700
rect 6657 -726 6687 -700
rect 6753 -731 6783 -700
rect 6849 -726 6879 -700
rect 6945 -731 6975 -700
rect 7041 -726 7071 -700
rect 7137 -731 7167 -700
rect 7233 -726 7263 -700
rect 7329 -731 7359 -700
rect 7425 -726 7455 -700
rect 7521 -731 7551 -700
rect 7617 -726 7647 -700
rect 7713 -731 7743 -700
rect 7809 -726 7839 -700
rect 7905 -731 7935 -700
rect 8001 -726 8031 -700
rect 8097 -731 8127 -700
rect 8193 -726 8223 -700
rect 8289 -731 8319 -700
rect 8385 -726 8415 -700
rect 8481 -731 8511 -700
rect 8577 -726 8607 -700
rect 8673 -731 8703 -700
rect 8769 -726 8799 -700
rect 8865 -731 8895 -700
rect 8961 -726 8991 -700
rect 9057 -731 9087 -700
rect 9153 -726 9183 -700
rect 9249 -731 9279 -700
rect 9345 -726 9375 -700
rect 9441 -731 9471 -700
rect 9537 -726 9567 -700
rect 9633 -731 9663 -700
rect 9729 -726 9759 -700
rect 9825 -731 9855 -700
rect 9921 -726 9951 -700
rect 10017 -731 10047 -700
rect 10113 -726 10143 -700
rect 10209 -731 10239 -700
rect 10305 -726 10335 -700
rect 10401 -731 10431 -700
rect 10497 -726 10527 -700
rect -10545 -747 -10479 -731
rect -10545 -781 -10529 -747
rect -10495 -781 -10479 -747
rect -10545 -797 -10479 -781
rect -10353 -747 -10287 -731
rect -10353 -781 -10337 -747
rect -10303 -781 -10287 -747
rect -10353 -797 -10287 -781
rect -10161 -747 -10095 -731
rect -10161 -781 -10145 -747
rect -10111 -781 -10095 -747
rect -10161 -797 -10095 -781
rect -9969 -747 -9903 -731
rect -9969 -781 -9953 -747
rect -9919 -781 -9903 -747
rect -9969 -797 -9903 -781
rect -9777 -747 -9711 -731
rect -9777 -781 -9761 -747
rect -9727 -781 -9711 -747
rect -9777 -797 -9711 -781
rect -9585 -747 -9519 -731
rect -9585 -781 -9569 -747
rect -9535 -781 -9519 -747
rect -9585 -797 -9519 -781
rect -9393 -747 -9327 -731
rect -9393 -781 -9377 -747
rect -9343 -781 -9327 -747
rect -9393 -797 -9327 -781
rect -9201 -747 -9135 -731
rect -9201 -781 -9185 -747
rect -9151 -781 -9135 -747
rect -9201 -797 -9135 -781
rect -9009 -747 -8943 -731
rect -9009 -781 -8993 -747
rect -8959 -781 -8943 -747
rect -9009 -797 -8943 -781
rect -8817 -747 -8751 -731
rect -8817 -781 -8801 -747
rect -8767 -781 -8751 -747
rect -8817 -797 -8751 -781
rect -8625 -747 -8559 -731
rect -8625 -781 -8609 -747
rect -8575 -781 -8559 -747
rect -8625 -797 -8559 -781
rect -8433 -747 -8367 -731
rect -8433 -781 -8417 -747
rect -8383 -781 -8367 -747
rect -8433 -797 -8367 -781
rect -8241 -747 -8175 -731
rect -8241 -781 -8225 -747
rect -8191 -781 -8175 -747
rect -8241 -797 -8175 -781
rect -8049 -747 -7983 -731
rect -8049 -781 -8033 -747
rect -7999 -781 -7983 -747
rect -8049 -797 -7983 -781
rect -7857 -747 -7791 -731
rect -7857 -781 -7841 -747
rect -7807 -781 -7791 -747
rect -7857 -797 -7791 -781
rect -7665 -747 -7599 -731
rect -7665 -781 -7649 -747
rect -7615 -781 -7599 -747
rect -7665 -797 -7599 -781
rect -7473 -747 -7407 -731
rect -7473 -781 -7457 -747
rect -7423 -781 -7407 -747
rect -7473 -797 -7407 -781
rect -7281 -747 -7215 -731
rect -7281 -781 -7265 -747
rect -7231 -781 -7215 -747
rect -7281 -797 -7215 -781
rect -7089 -747 -7023 -731
rect -7089 -781 -7073 -747
rect -7039 -781 -7023 -747
rect -7089 -797 -7023 -781
rect -6897 -747 -6831 -731
rect -6897 -781 -6881 -747
rect -6847 -781 -6831 -747
rect -6897 -797 -6831 -781
rect -6705 -747 -6639 -731
rect -6705 -781 -6689 -747
rect -6655 -781 -6639 -747
rect -6705 -797 -6639 -781
rect -6513 -747 -6447 -731
rect -6513 -781 -6497 -747
rect -6463 -781 -6447 -747
rect -6513 -797 -6447 -781
rect -6321 -747 -6255 -731
rect -6321 -781 -6305 -747
rect -6271 -781 -6255 -747
rect -6321 -797 -6255 -781
rect -6129 -747 -6063 -731
rect -6129 -781 -6113 -747
rect -6079 -781 -6063 -747
rect -6129 -797 -6063 -781
rect -5937 -747 -5871 -731
rect -5937 -781 -5921 -747
rect -5887 -781 -5871 -747
rect -5937 -797 -5871 -781
rect -5745 -747 -5679 -731
rect -5745 -781 -5729 -747
rect -5695 -781 -5679 -747
rect -5745 -797 -5679 -781
rect -5553 -747 -5487 -731
rect -5553 -781 -5537 -747
rect -5503 -781 -5487 -747
rect -5553 -797 -5487 -781
rect -5361 -747 -5295 -731
rect -5361 -781 -5345 -747
rect -5311 -781 -5295 -747
rect -5361 -797 -5295 -781
rect -5169 -747 -5103 -731
rect -5169 -781 -5153 -747
rect -5119 -781 -5103 -747
rect -5169 -797 -5103 -781
rect -4977 -747 -4911 -731
rect -4977 -781 -4961 -747
rect -4927 -781 -4911 -747
rect -4977 -797 -4911 -781
rect -4785 -747 -4719 -731
rect -4785 -781 -4769 -747
rect -4735 -781 -4719 -747
rect -4785 -797 -4719 -781
rect -4593 -747 -4527 -731
rect -4593 -781 -4577 -747
rect -4543 -781 -4527 -747
rect -4593 -797 -4527 -781
rect -4401 -747 -4335 -731
rect -4401 -781 -4385 -747
rect -4351 -781 -4335 -747
rect -4401 -797 -4335 -781
rect -4209 -747 -4143 -731
rect -4209 -781 -4193 -747
rect -4159 -781 -4143 -747
rect -4209 -797 -4143 -781
rect -4017 -747 -3951 -731
rect -4017 -781 -4001 -747
rect -3967 -781 -3951 -747
rect -4017 -797 -3951 -781
rect -3825 -747 -3759 -731
rect -3825 -781 -3809 -747
rect -3775 -781 -3759 -747
rect -3825 -797 -3759 -781
rect -3633 -747 -3567 -731
rect -3633 -781 -3617 -747
rect -3583 -781 -3567 -747
rect -3633 -797 -3567 -781
rect -3441 -747 -3375 -731
rect -3441 -781 -3425 -747
rect -3391 -781 -3375 -747
rect -3441 -797 -3375 -781
rect -3249 -747 -3183 -731
rect -3249 -781 -3233 -747
rect -3199 -781 -3183 -747
rect -3249 -797 -3183 -781
rect -3057 -747 -2991 -731
rect -3057 -781 -3041 -747
rect -3007 -781 -2991 -747
rect -3057 -797 -2991 -781
rect -2865 -747 -2799 -731
rect -2865 -781 -2849 -747
rect -2815 -781 -2799 -747
rect -2865 -797 -2799 -781
rect -2673 -747 -2607 -731
rect -2673 -781 -2657 -747
rect -2623 -781 -2607 -747
rect -2673 -797 -2607 -781
rect -2481 -747 -2415 -731
rect -2481 -781 -2465 -747
rect -2431 -781 -2415 -747
rect -2481 -797 -2415 -781
rect -2289 -747 -2223 -731
rect -2289 -781 -2273 -747
rect -2239 -781 -2223 -747
rect -2289 -797 -2223 -781
rect -2097 -747 -2031 -731
rect -2097 -781 -2081 -747
rect -2047 -781 -2031 -747
rect -2097 -797 -2031 -781
rect -1905 -747 -1839 -731
rect -1905 -781 -1889 -747
rect -1855 -781 -1839 -747
rect -1905 -797 -1839 -781
rect -1713 -747 -1647 -731
rect -1713 -781 -1697 -747
rect -1663 -781 -1647 -747
rect -1713 -797 -1647 -781
rect -1521 -747 -1455 -731
rect -1521 -781 -1505 -747
rect -1471 -781 -1455 -747
rect -1521 -797 -1455 -781
rect -1329 -747 -1263 -731
rect -1329 -781 -1313 -747
rect -1279 -781 -1263 -747
rect -1329 -797 -1263 -781
rect -1137 -747 -1071 -731
rect -1137 -781 -1121 -747
rect -1087 -781 -1071 -747
rect -1137 -797 -1071 -781
rect -945 -747 -879 -731
rect -945 -781 -929 -747
rect -895 -781 -879 -747
rect -945 -797 -879 -781
rect -753 -747 -687 -731
rect -753 -781 -737 -747
rect -703 -781 -687 -747
rect -753 -797 -687 -781
rect -561 -747 -495 -731
rect -561 -781 -545 -747
rect -511 -781 -495 -747
rect -561 -797 -495 -781
rect -369 -747 -303 -731
rect -369 -781 -353 -747
rect -319 -781 -303 -747
rect -369 -797 -303 -781
rect -177 -747 -111 -731
rect -177 -781 -161 -747
rect -127 -781 -111 -747
rect -177 -797 -111 -781
rect 15 -747 81 -731
rect 15 -781 31 -747
rect 65 -781 81 -747
rect 15 -797 81 -781
rect 207 -747 273 -731
rect 207 -781 223 -747
rect 257 -781 273 -747
rect 207 -797 273 -781
rect 399 -747 465 -731
rect 399 -781 415 -747
rect 449 -781 465 -747
rect 399 -797 465 -781
rect 591 -747 657 -731
rect 591 -781 607 -747
rect 641 -781 657 -747
rect 591 -797 657 -781
rect 783 -747 849 -731
rect 783 -781 799 -747
rect 833 -781 849 -747
rect 783 -797 849 -781
rect 975 -747 1041 -731
rect 975 -781 991 -747
rect 1025 -781 1041 -747
rect 975 -797 1041 -781
rect 1167 -747 1233 -731
rect 1167 -781 1183 -747
rect 1217 -781 1233 -747
rect 1167 -797 1233 -781
rect 1359 -747 1425 -731
rect 1359 -781 1375 -747
rect 1409 -781 1425 -747
rect 1359 -797 1425 -781
rect 1551 -747 1617 -731
rect 1551 -781 1567 -747
rect 1601 -781 1617 -747
rect 1551 -797 1617 -781
rect 1743 -747 1809 -731
rect 1743 -781 1759 -747
rect 1793 -781 1809 -747
rect 1743 -797 1809 -781
rect 1935 -747 2001 -731
rect 1935 -781 1951 -747
rect 1985 -781 2001 -747
rect 1935 -797 2001 -781
rect 2127 -747 2193 -731
rect 2127 -781 2143 -747
rect 2177 -781 2193 -747
rect 2127 -797 2193 -781
rect 2319 -747 2385 -731
rect 2319 -781 2335 -747
rect 2369 -781 2385 -747
rect 2319 -797 2385 -781
rect 2511 -747 2577 -731
rect 2511 -781 2527 -747
rect 2561 -781 2577 -747
rect 2511 -797 2577 -781
rect 2703 -747 2769 -731
rect 2703 -781 2719 -747
rect 2753 -781 2769 -747
rect 2703 -797 2769 -781
rect 2895 -747 2961 -731
rect 2895 -781 2911 -747
rect 2945 -781 2961 -747
rect 2895 -797 2961 -781
rect 3087 -747 3153 -731
rect 3087 -781 3103 -747
rect 3137 -781 3153 -747
rect 3087 -797 3153 -781
rect 3279 -747 3345 -731
rect 3279 -781 3295 -747
rect 3329 -781 3345 -747
rect 3279 -797 3345 -781
rect 3471 -747 3537 -731
rect 3471 -781 3487 -747
rect 3521 -781 3537 -747
rect 3471 -797 3537 -781
rect 3663 -747 3729 -731
rect 3663 -781 3679 -747
rect 3713 -781 3729 -747
rect 3663 -797 3729 -781
rect 3855 -747 3921 -731
rect 3855 -781 3871 -747
rect 3905 -781 3921 -747
rect 3855 -797 3921 -781
rect 4047 -747 4113 -731
rect 4047 -781 4063 -747
rect 4097 -781 4113 -747
rect 4047 -797 4113 -781
rect 4239 -747 4305 -731
rect 4239 -781 4255 -747
rect 4289 -781 4305 -747
rect 4239 -797 4305 -781
rect 4431 -747 4497 -731
rect 4431 -781 4447 -747
rect 4481 -781 4497 -747
rect 4431 -797 4497 -781
rect 4623 -747 4689 -731
rect 4623 -781 4639 -747
rect 4673 -781 4689 -747
rect 4623 -797 4689 -781
rect 4815 -747 4881 -731
rect 4815 -781 4831 -747
rect 4865 -781 4881 -747
rect 4815 -797 4881 -781
rect 5007 -747 5073 -731
rect 5007 -781 5023 -747
rect 5057 -781 5073 -747
rect 5007 -797 5073 -781
rect 5199 -747 5265 -731
rect 5199 -781 5215 -747
rect 5249 -781 5265 -747
rect 5199 -797 5265 -781
rect 5391 -747 5457 -731
rect 5391 -781 5407 -747
rect 5441 -781 5457 -747
rect 5391 -797 5457 -781
rect 5583 -747 5649 -731
rect 5583 -781 5599 -747
rect 5633 -781 5649 -747
rect 5583 -797 5649 -781
rect 5775 -747 5841 -731
rect 5775 -781 5791 -747
rect 5825 -781 5841 -747
rect 5775 -797 5841 -781
rect 5967 -747 6033 -731
rect 5967 -781 5983 -747
rect 6017 -781 6033 -747
rect 5967 -797 6033 -781
rect 6159 -747 6225 -731
rect 6159 -781 6175 -747
rect 6209 -781 6225 -747
rect 6159 -797 6225 -781
rect 6351 -747 6417 -731
rect 6351 -781 6367 -747
rect 6401 -781 6417 -747
rect 6351 -797 6417 -781
rect 6543 -747 6609 -731
rect 6543 -781 6559 -747
rect 6593 -781 6609 -747
rect 6543 -797 6609 -781
rect 6735 -747 6801 -731
rect 6735 -781 6751 -747
rect 6785 -781 6801 -747
rect 6735 -797 6801 -781
rect 6927 -747 6993 -731
rect 6927 -781 6943 -747
rect 6977 -781 6993 -747
rect 6927 -797 6993 -781
rect 7119 -747 7185 -731
rect 7119 -781 7135 -747
rect 7169 -781 7185 -747
rect 7119 -797 7185 -781
rect 7311 -747 7377 -731
rect 7311 -781 7327 -747
rect 7361 -781 7377 -747
rect 7311 -797 7377 -781
rect 7503 -747 7569 -731
rect 7503 -781 7519 -747
rect 7553 -781 7569 -747
rect 7503 -797 7569 -781
rect 7695 -747 7761 -731
rect 7695 -781 7711 -747
rect 7745 -781 7761 -747
rect 7695 -797 7761 -781
rect 7887 -747 7953 -731
rect 7887 -781 7903 -747
rect 7937 -781 7953 -747
rect 7887 -797 7953 -781
rect 8079 -747 8145 -731
rect 8079 -781 8095 -747
rect 8129 -781 8145 -747
rect 8079 -797 8145 -781
rect 8271 -747 8337 -731
rect 8271 -781 8287 -747
rect 8321 -781 8337 -747
rect 8271 -797 8337 -781
rect 8463 -747 8529 -731
rect 8463 -781 8479 -747
rect 8513 -781 8529 -747
rect 8463 -797 8529 -781
rect 8655 -747 8721 -731
rect 8655 -781 8671 -747
rect 8705 -781 8721 -747
rect 8655 -797 8721 -781
rect 8847 -747 8913 -731
rect 8847 -781 8863 -747
rect 8897 -781 8913 -747
rect 8847 -797 8913 -781
rect 9039 -747 9105 -731
rect 9039 -781 9055 -747
rect 9089 -781 9105 -747
rect 9039 -797 9105 -781
rect 9231 -747 9297 -731
rect 9231 -781 9247 -747
rect 9281 -781 9297 -747
rect 9231 -797 9297 -781
rect 9423 -747 9489 -731
rect 9423 -781 9439 -747
rect 9473 -781 9489 -747
rect 9423 -797 9489 -781
rect 9615 -747 9681 -731
rect 9615 -781 9631 -747
rect 9665 -781 9681 -747
rect 9615 -797 9681 -781
rect 9807 -747 9873 -731
rect 9807 -781 9823 -747
rect 9857 -781 9873 -747
rect 9807 -797 9873 -781
rect 9999 -747 10065 -731
rect 9999 -781 10015 -747
rect 10049 -781 10065 -747
rect 9999 -797 10065 -781
rect 10191 -747 10257 -731
rect 10191 -781 10207 -747
rect 10241 -781 10257 -747
rect 10191 -797 10257 -781
rect 10383 -747 10449 -731
rect 10383 -781 10399 -747
rect 10433 -781 10449 -747
rect 10383 -797 10449 -781
<< polycont >>
rect -10433 747 -10399 781
rect -10241 747 -10207 781
rect -10049 747 -10015 781
rect -9857 747 -9823 781
rect -9665 747 -9631 781
rect -9473 747 -9439 781
rect -9281 747 -9247 781
rect -9089 747 -9055 781
rect -8897 747 -8863 781
rect -8705 747 -8671 781
rect -8513 747 -8479 781
rect -8321 747 -8287 781
rect -8129 747 -8095 781
rect -7937 747 -7903 781
rect -7745 747 -7711 781
rect -7553 747 -7519 781
rect -7361 747 -7327 781
rect -7169 747 -7135 781
rect -6977 747 -6943 781
rect -6785 747 -6751 781
rect -6593 747 -6559 781
rect -6401 747 -6367 781
rect -6209 747 -6175 781
rect -6017 747 -5983 781
rect -5825 747 -5791 781
rect -5633 747 -5599 781
rect -5441 747 -5407 781
rect -5249 747 -5215 781
rect -5057 747 -5023 781
rect -4865 747 -4831 781
rect -4673 747 -4639 781
rect -4481 747 -4447 781
rect -4289 747 -4255 781
rect -4097 747 -4063 781
rect -3905 747 -3871 781
rect -3713 747 -3679 781
rect -3521 747 -3487 781
rect -3329 747 -3295 781
rect -3137 747 -3103 781
rect -2945 747 -2911 781
rect -2753 747 -2719 781
rect -2561 747 -2527 781
rect -2369 747 -2335 781
rect -2177 747 -2143 781
rect -1985 747 -1951 781
rect -1793 747 -1759 781
rect -1601 747 -1567 781
rect -1409 747 -1375 781
rect -1217 747 -1183 781
rect -1025 747 -991 781
rect -833 747 -799 781
rect -641 747 -607 781
rect -449 747 -415 781
rect -257 747 -223 781
rect -65 747 -31 781
rect 127 747 161 781
rect 319 747 353 781
rect 511 747 545 781
rect 703 747 737 781
rect 895 747 929 781
rect 1087 747 1121 781
rect 1279 747 1313 781
rect 1471 747 1505 781
rect 1663 747 1697 781
rect 1855 747 1889 781
rect 2047 747 2081 781
rect 2239 747 2273 781
rect 2431 747 2465 781
rect 2623 747 2657 781
rect 2815 747 2849 781
rect 3007 747 3041 781
rect 3199 747 3233 781
rect 3391 747 3425 781
rect 3583 747 3617 781
rect 3775 747 3809 781
rect 3967 747 4001 781
rect 4159 747 4193 781
rect 4351 747 4385 781
rect 4543 747 4577 781
rect 4735 747 4769 781
rect 4927 747 4961 781
rect 5119 747 5153 781
rect 5311 747 5345 781
rect 5503 747 5537 781
rect 5695 747 5729 781
rect 5887 747 5921 781
rect 6079 747 6113 781
rect 6271 747 6305 781
rect 6463 747 6497 781
rect 6655 747 6689 781
rect 6847 747 6881 781
rect 7039 747 7073 781
rect 7231 747 7265 781
rect 7423 747 7457 781
rect 7615 747 7649 781
rect 7807 747 7841 781
rect 7999 747 8033 781
rect 8191 747 8225 781
rect 8383 747 8417 781
rect 8575 747 8609 781
rect 8767 747 8801 781
rect 8959 747 8993 781
rect 9151 747 9185 781
rect 9343 747 9377 781
rect 9535 747 9569 781
rect 9727 747 9761 781
rect 9919 747 9953 781
rect 10111 747 10145 781
rect 10303 747 10337 781
rect 10495 747 10529 781
rect -10529 -781 -10495 -747
rect -10337 -781 -10303 -747
rect -10145 -781 -10111 -747
rect -9953 -781 -9919 -747
rect -9761 -781 -9727 -747
rect -9569 -781 -9535 -747
rect -9377 -781 -9343 -747
rect -9185 -781 -9151 -747
rect -8993 -781 -8959 -747
rect -8801 -781 -8767 -747
rect -8609 -781 -8575 -747
rect -8417 -781 -8383 -747
rect -8225 -781 -8191 -747
rect -8033 -781 -7999 -747
rect -7841 -781 -7807 -747
rect -7649 -781 -7615 -747
rect -7457 -781 -7423 -747
rect -7265 -781 -7231 -747
rect -7073 -781 -7039 -747
rect -6881 -781 -6847 -747
rect -6689 -781 -6655 -747
rect -6497 -781 -6463 -747
rect -6305 -781 -6271 -747
rect -6113 -781 -6079 -747
rect -5921 -781 -5887 -747
rect -5729 -781 -5695 -747
rect -5537 -781 -5503 -747
rect -5345 -781 -5311 -747
rect -5153 -781 -5119 -747
rect -4961 -781 -4927 -747
rect -4769 -781 -4735 -747
rect -4577 -781 -4543 -747
rect -4385 -781 -4351 -747
rect -4193 -781 -4159 -747
rect -4001 -781 -3967 -747
rect -3809 -781 -3775 -747
rect -3617 -781 -3583 -747
rect -3425 -781 -3391 -747
rect -3233 -781 -3199 -747
rect -3041 -781 -3007 -747
rect -2849 -781 -2815 -747
rect -2657 -781 -2623 -747
rect -2465 -781 -2431 -747
rect -2273 -781 -2239 -747
rect -2081 -781 -2047 -747
rect -1889 -781 -1855 -747
rect -1697 -781 -1663 -747
rect -1505 -781 -1471 -747
rect -1313 -781 -1279 -747
rect -1121 -781 -1087 -747
rect -929 -781 -895 -747
rect -737 -781 -703 -747
rect -545 -781 -511 -747
rect -353 -781 -319 -747
rect -161 -781 -127 -747
rect 31 -781 65 -747
rect 223 -781 257 -747
rect 415 -781 449 -747
rect 607 -781 641 -747
rect 799 -781 833 -747
rect 991 -781 1025 -747
rect 1183 -781 1217 -747
rect 1375 -781 1409 -747
rect 1567 -781 1601 -747
rect 1759 -781 1793 -747
rect 1951 -781 1985 -747
rect 2143 -781 2177 -747
rect 2335 -781 2369 -747
rect 2527 -781 2561 -747
rect 2719 -781 2753 -747
rect 2911 -781 2945 -747
rect 3103 -781 3137 -747
rect 3295 -781 3329 -747
rect 3487 -781 3521 -747
rect 3679 -781 3713 -747
rect 3871 -781 3905 -747
rect 4063 -781 4097 -747
rect 4255 -781 4289 -747
rect 4447 -781 4481 -747
rect 4639 -781 4673 -747
rect 4831 -781 4865 -747
rect 5023 -781 5057 -747
rect 5215 -781 5249 -747
rect 5407 -781 5441 -747
rect 5599 -781 5633 -747
rect 5791 -781 5825 -747
rect 5983 -781 6017 -747
rect 6175 -781 6209 -747
rect 6367 -781 6401 -747
rect 6559 -781 6593 -747
rect 6751 -781 6785 -747
rect 6943 -781 6977 -747
rect 7135 -781 7169 -747
rect 7327 -781 7361 -747
rect 7519 -781 7553 -747
rect 7711 -781 7745 -747
rect 7903 -781 7937 -747
rect 8095 -781 8129 -747
rect 8287 -781 8321 -747
rect 8479 -781 8513 -747
rect 8671 -781 8705 -747
rect 8863 -781 8897 -747
rect 9055 -781 9089 -747
rect 9247 -781 9281 -747
rect 9439 -781 9473 -747
rect 9631 -781 9665 -747
rect 9823 -781 9857 -747
rect 10015 -781 10049 -747
rect 10207 -781 10241 -747
rect 10399 -781 10433 -747
<< locali >>
rect -10691 849 -10595 883
rect 10595 849 10691 883
rect -10691 787 -10657 849
rect 10657 787 10691 849
rect -10449 747 -10433 781
rect -10399 747 -10383 781
rect -10257 747 -10241 781
rect -10207 747 -10191 781
rect -10065 747 -10049 781
rect -10015 747 -9999 781
rect -9873 747 -9857 781
rect -9823 747 -9807 781
rect -9681 747 -9665 781
rect -9631 747 -9615 781
rect -9489 747 -9473 781
rect -9439 747 -9423 781
rect -9297 747 -9281 781
rect -9247 747 -9231 781
rect -9105 747 -9089 781
rect -9055 747 -9039 781
rect -8913 747 -8897 781
rect -8863 747 -8847 781
rect -8721 747 -8705 781
rect -8671 747 -8655 781
rect -8529 747 -8513 781
rect -8479 747 -8463 781
rect -8337 747 -8321 781
rect -8287 747 -8271 781
rect -8145 747 -8129 781
rect -8095 747 -8079 781
rect -7953 747 -7937 781
rect -7903 747 -7887 781
rect -7761 747 -7745 781
rect -7711 747 -7695 781
rect -7569 747 -7553 781
rect -7519 747 -7503 781
rect -7377 747 -7361 781
rect -7327 747 -7311 781
rect -7185 747 -7169 781
rect -7135 747 -7119 781
rect -6993 747 -6977 781
rect -6943 747 -6927 781
rect -6801 747 -6785 781
rect -6751 747 -6735 781
rect -6609 747 -6593 781
rect -6559 747 -6543 781
rect -6417 747 -6401 781
rect -6367 747 -6351 781
rect -6225 747 -6209 781
rect -6175 747 -6159 781
rect -6033 747 -6017 781
rect -5983 747 -5967 781
rect -5841 747 -5825 781
rect -5791 747 -5775 781
rect -5649 747 -5633 781
rect -5599 747 -5583 781
rect -5457 747 -5441 781
rect -5407 747 -5391 781
rect -5265 747 -5249 781
rect -5215 747 -5199 781
rect -5073 747 -5057 781
rect -5023 747 -5007 781
rect -4881 747 -4865 781
rect -4831 747 -4815 781
rect -4689 747 -4673 781
rect -4639 747 -4623 781
rect -4497 747 -4481 781
rect -4447 747 -4431 781
rect -4305 747 -4289 781
rect -4255 747 -4239 781
rect -4113 747 -4097 781
rect -4063 747 -4047 781
rect -3921 747 -3905 781
rect -3871 747 -3855 781
rect -3729 747 -3713 781
rect -3679 747 -3663 781
rect -3537 747 -3521 781
rect -3487 747 -3471 781
rect -3345 747 -3329 781
rect -3295 747 -3279 781
rect -3153 747 -3137 781
rect -3103 747 -3087 781
rect -2961 747 -2945 781
rect -2911 747 -2895 781
rect -2769 747 -2753 781
rect -2719 747 -2703 781
rect -2577 747 -2561 781
rect -2527 747 -2511 781
rect -2385 747 -2369 781
rect -2335 747 -2319 781
rect -2193 747 -2177 781
rect -2143 747 -2127 781
rect -2001 747 -1985 781
rect -1951 747 -1935 781
rect -1809 747 -1793 781
rect -1759 747 -1743 781
rect -1617 747 -1601 781
rect -1567 747 -1551 781
rect -1425 747 -1409 781
rect -1375 747 -1359 781
rect -1233 747 -1217 781
rect -1183 747 -1167 781
rect -1041 747 -1025 781
rect -991 747 -975 781
rect -849 747 -833 781
rect -799 747 -783 781
rect -657 747 -641 781
rect -607 747 -591 781
rect -465 747 -449 781
rect -415 747 -399 781
rect -273 747 -257 781
rect -223 747 -207 781
rect -81 747 -65 781
rect -31 747 -15 781
rect 111 747 127 781
rect 161 747 177 781
rect 303 747 319 781
rect 353 747 369 781
rect 495 747 511 781
rect 545 747 561 781
rect 687 747 703 781
rect 737 747 753 781
rect 879 747 895 781
rect 929 747 945 781
rect 1071 747 1087 781
rect 1121 747 1137 781
rect 1263 747 1279 781
rect 1313 747 1329 781
rect 1455 747 1471 781
rect 1505 747 1521 781
rect 1647 747 1663 781
rect 1697 747 1713 781
rect 1839 747 1855 781
rect 1889 747 1905 781
rect 2031 747 2047 781
rect 2081 747 2097 781
rect 2223 747 2239 781
rect 2273 747 2289 781
rect 2415 747 2431 781
rect 2465 747 2481 781
rect 2607 747 2623 781
rect 2657 747 2673 781
rect 2799 747 2815 781
rect 2849 747 2865 781
rect 2991 747 3007 781
rect 3041 747 3057 781
rect 3183 747 3199 781
rect 3233 747 3249 781
rect 3375 747 3391 781
rect 3425 747 3441 781
rect 3567 747 3583 781
rect 3617 747 3633 781
rect 3759 747 3775 781
rect 3809 747 3825 781
rect 3951 747 3967 781
rect 4001 747 4017 781
rect 4143 747 4159 781
rect 4193 747 4209 781
rect 4335 747 4351 781
rect 4385 747 4401 781
rect 4527 747 4543 781
rect 4577 747 4593 781
rect 4719 747 4735 781
rect 4769 747 4785 781
rect 4911 747 4927 781
rect 4961 747 4977 781
rect 5103 747 5119 781
rect 5153 747 5169 781
rect 5295 747 5311 781
rect 5345 747 5361 781
rect 5487 747 5503 781
rect 5537 747 5553 781
rect 5679 747 5695 781
rect 5729 747 5745 781
rect 5871 747 5887 781
rect 5921 747 5937 781
rect 6063 747 6079 781
rect 6113 747 6129 781
rect 6255 747 6271 781
rect 6305 747 6321 781
rect 6447 747 6463 781
rect 6497 747 6513 781
rect 6639 747 6655 781
rect 6689 747 6705 781
rect 6831 747 6847 781
rect 6881 747 6897 781
rect 7023 747 7039 781
rect 7073 747 7089 781
rect 7215 747 7231 781
rect 7265 747 7281 781
rect 7407 747 7423 781
rect 7457 747 7473 781
rect 7599 747 7615 781
rect 7649 747 7665 781
rect 7791 747 7807 781
rect 7841 747 7857 781
rect 7983 747 7999 781
rect 8033 747 8049 781
rect 8175 747 8191 781
rect 8225 747 8241 781
rect 8367 747 8383 781
rect 8417 747 8433 781
rect 8559 747 8575 781
rect 8609 747 8625 781
rect 8751 747 8767 781
rect 8801 747 8817 781
rect 8943 747 8959 781
rect 8993 747 9009 781
rect 9135 747 9151 781
rect 9185 747 9201 781
rect 9327 747 9343 781
rect 9377 747 9393 781
rect 9519 747 9535 781
rect 9569 747 9585 781
rect 9711 747 9727 781
rect 9761 747 9777 781
rect 9903 747 9919 781
rect 9953 747 9969 781
rect 10095 747 10111 781
rect 10145 747 10161 781
rect 10287 747 10303 781
rect 10337 747 10353 781
rect 10479 747 10495 781
rect 10529 747 10545 781
rect -10577 688 -10543 704
rect -10577 -704 -10543 -688
rect -10481 688 -10447 704
rect -10481 -704 -10447 -688
rect -10385 688 -10351 704
rect -10385 -704 -10351 -688
rect -10289 688 -10255 704
rect -10289 -704 -10255 -688
rect -10193 688 -10159 704
rect -10193 -704 -10159 -688
rect -10097 688 -10063 704
rect -10097 -704 -10063 -688
rect -10001 688 -9967 704
rect -10001 -704 -9967 -688
rect -9905 688 -9871 704
rect -9905 -704 -9871 -688
rect -9809 688 -9775 704
rect -9809 -704 -9775 -688
rect -9713 688 -9679 704
rect -9713 -704 -9679 -688
rect -9617 688 -9583 704
rect -9617 -704 -9583 -688
rect -9521 688 -9487 704
rect -9521 -704 -9487 -688
rect -9425 688 -9391 704
rect -9425 -704 -9391 -688
rect -9329 688 -9295 704
rect -9329 -704 -9295 -688
rect -9233 688 -9199 704
rect -9233 -704 -9199 -688
rect -9137 688 -9103 704
rect -9137 -704 -9103 -688
rect -9041 688 -9007 704
rect -9041 -704 -9007 -688
rect -8945 688 -8911 704
rect -8945 -704 -8911 -688
rect -8849 688 -8815 704
rect -8849 -704 -8815 -688
rect -8753 688 -8719 704
rect -8753 -704 -8719 -688
rect -8657 688 -8623 704
rect -8657 -704 -8623 -688
rect -8561 688 -8527 704
rect -8561 -704 -8527 -688
rect -8465 688 -8431 704
rect -8465 -704 -8431 -688
rect -8369 688 -8335 704
rect -8369 -704 -8335 -688
rect -8273 688 -8239 704
rect -8273 -704 -8239 -688
rect -8177 688 -8143 704
rect -8177 -704 -8143 -688
rect -8081 688 -8047 704
rect -8081 -704 -8047 -688
rect -7985 688 -7951 704
rect -7985 -704 -7951 -688
rect -7889 688 -7855 704
rect -7889 -704 -7855 -688
rect -7793 688 -7759 704
rect -7793 -704 -7759 -688
rect -7697 688 -7663 704
rect -7697 -704 -7663 -688
rect -7601 688 -7567 704
rect -7601 -704 -7567 -688
rect -7505 688 -7471 704
rect -7505 -704 -7471 -688
rect -7409 688 -7375 704
rect -7409 -704 -7375 -688
rect -7313 688 -7279 704
rect -7313 -704 -7279 -688
rect -7217 688 -7183 704
rect -7217 -704 -7183 -688
rect -7121 688 -7087 704
rect -7121 -704 -7087 -688
rect -7025 688 -6991 704
rect -7025 -704 -6991 -688
rect -6929 688 -6895 704
rect -6929 -704 -6895 -688
rect -6833 688 -6799 704
rect -6833 -704 -6799 -688
rect -6737 688 -6703 704
rect -6737 -704 -6703 -688
rect -6641 688 -6607 704
rect -6641 -704 -6607 -688
rect -6545 688 -6511 704
rect -6545 -704 -6511 -688
rect -6449 688 -6415 704
rect -6449 -704 -6415 -688
rect -6353 688 -6319 704
rect -6353 -704 -6319 -688
rect -6257 688 -6223 704
rect -6257 -704 -6223 -688
rect -6161 688 -6127 704
rect -6161 -704 -6127 -688
rect -6065 688 -6031 704
rect -6065 -704 -6031 -688
rect -5969 688 -5935 704
rect -5969 -704 -5935 -688
rect -5873 688 -5839 704
rect -5873 -704 -5839 -688
rect -5777 688 -5743 704
rect -5777 -704 -5743 -688
rect -5681 688 -5647 704
rect -5681 -704 -5647 -688
rect -5585 688 -5551 704
rect -5585 -704 -5551 -688
rect -5489 688 -5455 704
rect -5489 -704 -5455 -688
rect -5393 688 -5359 704
rect -5393 -704 -5359 -688
rect -5297 688 -5263 704
rect -5297 -704 -5263 -688
rect -5201 688 -5167 704
rect -5201 -704 -5167 -688
rect -5105 688 -5071 704
rect -5105 -704 -5071 -688
rect -5009 688 -4975 704
rect -5009 -704 -4975 -688
rect -4913 688 -4879 704
rect -4913 -704 -4879 -688
rect -4817 688 -4783 704
rect -4817 -704 -4783 -688
rect -4721 688 -4687 704
rect -4721 -704 -4687 -688
rect -4625 688 -4591 704
rect -4625 -704 -4591 -688
rect -4529 688 -4495 704
rect -4529 -704 -4495 -688
rect -4433 688 -4399 704
rect -4433 -704 -4399 -688
rect -4337 688 -4303 704
rect -4337 -704 -4303 -688
rect -4241 688 -4207 704
rect -4241 -704 -4207 -688
rect -4145 688 -4111 704
rect -4145 -704 -4111 -688
rect -4049 688 -4015 704
rect -4049 -704 -4015 -688
rect -3953 688 -3919 704
rect -3953 -704 -3919 -688
rect -3857 688 -3823 704
rect -3857 -704 -3823 -688
rect -3761 688 -3727 704
rect -3761 -704 -3727 -688
rect -3665 688 -3631 704
rect -3665 -704 -3631 -688
rect -3569 688 -3535 704
rect -3569 -704 -3535 -688
rect -3473 688 -3439 704
rect -3473 -704 -3439 -688
rect -3377 688 -3343 704
rect -3377 -704 -3343 -688
rect -3281 688 -3247 704
rect -3281 -704 -3247 -688
rect -3185 688 -3151 704
rect -3185 -704 -3151 -688
rect -3089 688 -3055 704
rect -3089 -704 -3055 -688
rect -2993 688 -2959 704
rect -2993 -704 -2959 -688
rect -2897 688 -2863 704
rect -2897 -704 -2863 -688
rect -2801 688 -2767 704
rect -2801 -704 -2767 -688
rect -2705 688 -2671 704
rect -2705 -704 -2671 -688
rect -2609 688 -2575 704
rect -2609 -704 -2575 -688
rect -2513 688 -2479 704
rect -2513 -704 -2479 -688
rect -2417 688 -2383 704
rect -2417 -704 -2383 -688
rect -2321 688 -2287 704
rect -2321 -704 -2287 -688
rect -2225 688 -2191 704
rect -2225 -704 -2191 -688
rect -2129 688 -2095 704
rect -2129 -704 -2095 -688
rect -2033 688 -1999 704
rect -2033 -704 -1999 -688
rect -1937 688 -1903 704
rect -1937 -704 -1903 -688
rect -1841 688 -1807 704
rect -1841 -704 -1807 -688
rect -1745 688 -1711 704
rect -1745 -704 -1711 -688
rect -1649 688 -1615 704
rect -1649 -704 -1615 -688
rect -1553 688 -1519 704
rect -1553 -704 -1519 -688
rect -1457 688 -1423 704
rect -1457 -704 -1423 -688
rect -1361 688 -1327 704
rect -1361 -704 -1327 -688
rect -1265 688 -1231 704
rect -1265 -704 -1231 -688
rect -1169 688 -1135 704
rect -1169 -704 -1135 -688
rect -1073 688 -1039 704
rect -1073 -704 -1039 -688
rect -977 688 -943 704
rect -977 -704 -943 -688
rect -881 688 -847 704
rect -881 -704 -847 -688
rect -785 688 -751 704
rect -785 -704 -751 -688
rect -689 688 -655 704
rect -689 -704 -655 -688
rect -593 688 -559 704
rect -593 -704 -559 -688
rect -497 688 -463 704
rect -497 -704 -463 -688
rect -401 688 -367 704
rect -401 -704 -367 -688
rect -305 688 -271 704
rect -305 -704 -271 -688
rect -209 688 -175 704
rect -209 -704 -175 -688
rect -113 688 -79 704
rect -113 -704 -79 -688
rect -17 688 17 704
rect -17 -704 17 -688
rect 79 688 113 704
rect 79 -704 113 -688
rect 175 688 209 704
rect 175 -704 209 -688
rect 271 688 305 704
rect 271 -704 305 -688
rect 367 688 401 704
rect 367 -704 401 -688
rect 463 688 497 704
rect 463 -704 497 -688
rect 559 688 593 704
rect 559 -704 593 -688
rect 655 688 689 704
rect 655 -704 689 -688
rect 751 688 785 704
rect 751 -704 785 -688
rect 847 688 881 704
rect 847 -704 881 -688
rect 943 688 977 704
rect 943 -704 977 -688
rect 1039 688 1073 704
rect 1039 -704 1073 -688
rect 1135 688 1169 704
rect 1135 -704 1169 -688
rect 1231 688 1265 704
rect 1231 -704 1265 -688
rect 1327 688 1361 704
rect 1327 -704 1361 -688
rect 1423 688 1457 704
rect 1423 -704 1457 -688
rect 1519 688 1553 704
rect 1519 -704 1553 -688
rect 1615 688 1649 704
rect 1615 -704 1649 -688
rect 1711 688 1745 704
rect 1711 -704 1745 -688
rect 1807 688 1841 704
rect 1807 -704 1841 -688
rect 1903 688 1937 704
rect 1903 -704 1937 -688
rect 1999 688 2033 704
rect 1999 -704 2033 -688
rect 2095 688 2129 704
rect 2095 -704 2129 -688
rect 2191 688 2225 704
rect 2191 -704 2225 -688
rect 2287 688 2321 704
rect 2287 -704 2321 -688
rect 2383 688 2417 704
rect 2383 -704 2417 -688
rect 2479 688 2513 704
rect 2479 -704 2513 -688
rect 2575 688 2609 704
rect 2575 -704 2609 -688
rect 2671 688 2705 704
rect 2671 -704 2705 -688
rect 2767 688 2801 704
rect 2767 -704 2801 -688
rect 2863 688 2897 704
rect 2863 -704 2897 -688
rect 2959 688 2993 704
rect 2959 -704 2993 -688
rect 3055 688 3089 704
rect 3055 -704 3089 -688
rect 3151 688 3185 704
rect 3151 -704 3185 -688
rect 3247 688 3281 704
rect 3247 -704 3281 -688
rect 3343 688 3377 704
rect 3343 -704 3377 -688
rect 3439 688 3473 704
rect 3439 -704 3473 -688
rect 3535 688 3569 704
rect 3535 -704 3569 -688
rect 3631 688 3665 704
rect 3631 -704 3665 -688
rect 3727 688 3761 704
rect 3727 -704 3761 -688
rect 3823 688 3857 704
rect 3823 -704 3857 -688
rect 3919 688 3953 704
rect 3919 -704 3953 -688
rect 4015 688 4049 704
rect 4015 -704 4049 -688
rect 4111 688 4145 704
rect 4111 -704 4145 -688
rect 4207 688 4241 704
rect 4207 -704 4241 -688
rect 4303 688 4337 704
rect 4303 -704 4337 -688
rect 4399 688 4433 704
rect 4399 -704 4433 -688
rect 4495 688 4529 704
rect 4495 -704 4529 -688
rect 4591 688 4625 704
rect 4591 -704 4625 -688
rect 4687 688 4721 704
rect 4687 -704 4721 -688
rect 4783 688 4817 704
rect 4783 -704 4817 -688
rect 4879 688 4913 704
rect 4879 -704 4913 -688
rect 4975 688 5009 704
rect 4975 -704 5009 -688
rect 5071 688 5105 704
rect 5071 -704 5105 -688
rect 5167 688 5201 704
rect 5167 -704 5201 -688
rect 5263 688 5297 704
rect 5263 -704 5297 -688
rect 5359 688 5393 704
rect 5359 -704 5393 -688
rect 5455 688 5489 704
rect 5455 -704 5489 -688
rect 5551 688 5585 704
rect 5551 -704 5585 -688
rect 5647 688 5681 704
rect 5647 -704 5681 -688
rect 5743 688 5777 704
rect 5743 -704 5777 -688
rect 5839 688 5873 704
rect 5839 -704 5873 -688
rect 5935 688 5969 704
rect 5935 -704 5969 -688
rect 6031 688 6065 704
rect 6031 -704 6065 -688
rect 6127 688 6161 704
rect 6127 -704 6161 -688
rect 6223 688 6257 704
rect 6223 -704 6257 -688
rect 6319 688 6353 704
rect 6319 -704 6353 -688
rect 6415 688 6449 704
rect 6415 -704 6449 -688
rect 6511 688 6545 704
rect 6511 -704 6545 -688
rect 6607 688 6641 704
rect 6607 -704 6641 -688
rect 6703 688 6737 704
rect 6703 -704 6737 -688
rect 6799 688 6833 704
rect 6799 -704 6833 -688
rect 6895 688 6929 704
rect 6895 -704 6929 -688
rect 6991 688 7025 704
rect 6991 -704 7025 -688
rect 7087 688 7121 704
rect 7087 -704 7121 -688
rect 7183 688 7217 704
rect 7183 -704 7217 -688
rect 7279 688 7313 704
rect 7279 -704 7313 -688
rect 7375 688 7409 704
rect 7375 -704 7409 -688
rect 7471 688 7505 704
rect 7471 -704 7505 -688
rect 7567 688 7601 704
rect 7567 -704 7601 -688
rect 7663 688 7697 704
rect 7663 -704 7697 -688
rect 7759 688 7793 704
rect 7759 -704 7793 -688
rect 7855 688 7889 704
rect 7855 -704 7889 -688
rect 7951 688 7985 704
rect 7951 -704 7985 -688
rect 8047 688 8081 704
rect 8047 -704 8081 -688
rect 8143 688 8177 704
rect 8143 -704 8177 -688
rect 8239 688 8273 704
rect 8239 -704 8273 -688
rect 8335 688 8369 704
rect 8335 -704 8369 -688
rect 8431 688 8465 704
rect 8431 -704 8465 -688
rect 8527 688 8561 704
rect 8527 -704 8561 -688
rect 8623 688 8657 704
rect 8623 -704 8657 -688
rect 8719 688 8753 704
rect 8719 -704 8753 -688
rect 8815 688 8849 704
rect 8815 -704 8849 -688
rect 8911 688 8945 704
rect 8911 -704 8945 -688
rect 9007 688 9041 704
rect 9007 -704 9041 -688
rect 9103 688 9137 704
rect 9103 -704 9137 -688
rect 9199 688 9233 704
rect 9199 -704 9233 -688
rect 9295 688 9329 704
rect 9295 -704 9329 -688
rect 9391 688 9425 704
rect 9391 -704 9425 -688
rect 9487 688 9521 704
rect 9487 -704 9521 -688
rect 9583 688 9617 704
rect 9583 -704 9617 -688
rect 9679 688 9713 704
rect 9679 -704 9713 -688
rect 9775 688 9809 704
rect 9775 -704 9809 -688
rect 9871 688 9905 704
rect 9871 -704 9905 -688
rect 9967 688 10001 704
rect 9967 -704 10001 -688
rect 10063 688 10097 704
rect 10063 -704 10097 -688
rect 10159 688 10193 704
rect 10159 -704 10193 -688
rect 10255 688 10289 704
rect 10255 -704 10289 -688
rect 10351 688 10385 704
rect 10351 -704 10385 -688
rect 10447 688 10481 704
rect 10447 -704 10481 -688
rect 10543 688 10577 704
rect 10543 -704 10577 -688
rect -10545 -781 -10529 -747
rect -10495 -781 -10479 -747
rect -10353 -781 -10337 -747
rect -10303 -781 -10287 -747
rect -10161 -781 -10145 -747
rect -10111 -781 -10095 -747
rect -9969 -781 -9953 -747
rect -9919 -781 -9903 -747
rect -9777 -781 -9761 -747
rect -9727 -781 -9711 -747
rect -9585 -781 -9569 -747
rect -9535 -781 -9519 -747
rect -9393 -781 -9377 -747
rect -9343 -781 -9327 -747
rect -9201 -781 -9185 -747
rect -9151 -781 -9135 -747
rect -9009 -781 -8993 -747
rect -8959 -781 -8943 -747
rect -8817 -781 -8801 -747
rect -8767 -781 -8751 -747
rect -8625 -781 -8609 -747
rect -8575 -781 -8559 -747
rect -8433 -781 -8417 -747
rect -8383 -781 -8367 -747
rect -8241 -781 -8225 -747
rect -8191 -781 -8175 -747
rect -8049 -781 -8033 -747
rect -7999 -781 -7983 -747
rect -7857 -781 -7841 -747
rect -7807 -781 -7791 -747
rect -7665 -781 -7649 -747
rect -7615 -781 -7599 -747
rect -7473 -781 -7457 -747
rect -7423 -781 -7407 -747
rect -7281 -781 -7265 -747
rect -7231 -781 -7215 -747
rect -7089 -781 -7073 -747
rect -7039 -781 -7023 -747
rect -6897 -781 -6881 -747
rect -6847 -781 -6831 -747
rect -6705 -781 -6689 -747
rect -6655 -781 -6639 -747
rect -6513 -781 -6497 -747
rect -6463 -781 -6447 -747
rect -6321 -781 -6305 -747
rect -6271 -781 -6255 -747
rect -6129 -781 -6113 -747
rect -6079 -781 -6063 -747
rect -5937 -781 -5921 -747
rect -5887 -781 -5871 -747
rect -5745 -781 -5729 -747
rect -5695 -781 -5679 -747
rect -5553 -781 -5537 -747
rect -5503 -781 -5487 -747
rect -5361 -781 -5345 -747
rect -5311 -781 -5295 -747
rect -5169 -781 -5153 -747
rect -5119 -781 -5103 -747
rect -4977 -781 -4961 -747
rect -4927 -781 -4911 -747
rect -4785 -781 -4769 -747
rect -4735 -781 -4719 -747
rect -4593 -781 -4577 -747
rect -4543 -781 -4527 -747
rect -4401 -781 -4385 -747
rect -4351 -781 -4335 -747
rect -4209 -781 -4193 -747
rect -4159 -781 -4143 -747
rect -4017 -781 -4001 -747
rect -3967 -781 -3951 -747
rect -3825 -781 -3809 -747
rect -3775 -781 -3759 -747
rect -3633 -781 -3617 -747
rect -3583 -781 -3567 -747
rect -3441 -781 -3425 -747
rect -3391 -781 -3375 -747
rect -3249 -781 -3233 -747
rect -3199 -781 -3183 -747
rect -3057 -781 -3041 -747
rect -3007 -781 -2991 -747
rect -2865 -781 -2849 -747
rect -2815 -781 -2799 -747
rect -2673 -781 -2657 -747
rect -2623 -781 -2607 -747
rect -2481 -781 -2465 -747
rect -2431 -781 -2415 -747
rect -2289 -781 -2273 -747
rect -2239 -781 -2223 -747
rect -2097 -781 -2081 -747
rect -2047 -781 -2031 -747
rect -1905 -781 -1889 -747
rect -1855 -781 -1839 -747
rect -1713 -781 -1697 -747
rect -1663 -781 -1647 -747
rect -1521 -781 -1505 -747
rect -1471 -781 -1455 -747
rect -1329 -781 -1313 -747
rect -1279 -781 -1263 -747
rect -1137 -781 -1121 -747
rect -1087 -781 -1071 -747
rect -945 -781 -929 -747
rect -895 -781 -879 -747
rect -753 -781 -737 -747
rect -703 -781 -687 -747
rect -561 -781 -545 -747
rect -511 -781 -495 -747
rect -369 -781 -353 -747
rect -319 -781 -303 -747
rect -177 -781 -161 -747
rect -127 -781 -111 -747
rect 15 -781 31 -747
rect 65 -781 81 -747
rect 207 -781 223 -747
rect 257 -781 273 -747
rect 399 -781 415 -747
rect 449 -781 465 -747
rect 591 -781 607 -747
rect 641 -781 657 -747
rect 783 -781 799 -747
rect 833 -781 849 -747
rect 975 -781 991 -747
rect 1025 -781 1041 -747
rect 1167 -781 1183 -747
rect 1217 -781 1233 -747
rect 1359 -781 1375 -747
rect 1409 -781 1425 -747
rect 1551 -781 1567 -747
rect 1601 -781 1617 -747
rect 1743 -781 1759 -747
rect 1793 -781 1809 -747
rect 1935 -781 1951 -747
rect 1985 -781 2001 -747
rect 2127 -781 2143 -747
rect 2177 -781 2193 -747
rect 2319 -781 2335 -747
rect 2369 -781 2385 -747
rect 2511 -781 2527 -747
rect 2561 -781 2577 -747
rect 2703 -781 2719 -747
rect 2753 -781 2769 -747
rect 2895 -781 2911 -747
rect 2945 -781 2961 -747
rect 3087 -781 3103 -747
rect 3137 -781 3153 -747
rect 3279 -781 3295 -747
rect 3329 -781 3345 -747
rect 3471 -781 3487 -747
rect 3521 -781 3537 -747
rect 3663 -781 3679 -747
rect 3713 -781 3729 -747
rect 3855 -781 3871 -747
rect 3905 -781 3921 -747
rect 4047 -781 4063 -747
rect 4097 -781 4113 -747
rect 4239 -781 4255 -747
rect 4289 -781 4305 -747
rect 4431 -781 4447 -747
rect 4481 -781 4497 -747
rect 4623 -781 4639 -747
rect 4673 -781 4689 -747
rect 4815 -781 4831 -747
rect 4865 -781 4881 -747
rect 5007 -781 5023 -747
rect 5057 -781 5073 -747
rect 5199 -781 5215 -747
rect 5249 -781 5265 -747
rect 5391 -781 5407 -747
rect 5441 -781 5457 -747
rect 5583 -781 5599 -747
rect 5633 -781 5649 -747
rect 5775 -781 5791 -747
rect 5825 -781 5841 -747
rect 5967 -781 5983 -747
rect 6017 -781 6033 -747
rect 6159 -781 6175 -747
rect 6209 -781 6225 -747
rect 6351 -781 6367 -747
rect 6401 -781 6417 -747
rect 6543 -781 6559 -747
rect 6593 -781 6609 -747
rect 6735 -781 6751 -747
rect 6785 -781 6801 -747
rect 6927 -781 6943 -747
rect 6977 -781 6993 -747
rect 7119 -781 7135 -747
rect 7169 -781 7185 -747
rect 7311 -781 7327 -747
rect 7361 -781 7377 -747
rect 7503 -781 7519 -747
rect 7553 -781 7569 -747
rect 7695 -781 7711 -747
rect 7745 -781 7761 -747
rect 7887 -781 7903 -747
rect 7937 -781 7953 -747
rect 8079 -781 8095 -747
rect 8129 -781 8145 -747
rect 8271 -781 8287 -747
rect 8321 -781 8337 -747
rect 8463 -781 8479 -747
rect 8513 -781 8529 -747
rect 8655 -781 8671 -747
rect 8705 -781 8721 -747
rect 8847 -781 8863 -747
rect 8897 -781 8913 -747
rect 9039 -781 9055 -747
rect 9089 -781 9105 -747
rect 9231 -781 9247 -747
rect 9281 -781 9297 -747
rect 9423 -781 9439 -747
rect 9473 -781 9489 -747
rect 9615 -781 9631 -747
rect 9665 -781 9681 -747
rect 9807 -781 9823 -747
rect 9857 -781 9873 -747
rect 9999 -781 10015 -747
rect 10049 -781 10065 -747
rect 10191 -781 10207 -747
rect 10241 -781 10257 -747
rect 10383 -781 10399 -747
rect 10433 -781 10449 -747
rect -10691 -849 -10657 -787
rect 10657 -849 10691 -787
rect -10691 -883 -10595 -849
rect 10595 -883 10691 -849
<< viali >>
rect -10433 747 -10399 781
rect -10241 747 -10207 781
rect -10049 747 -10015 781
rect -9857 747 -9823 781
rect -9665 747 -9631 781
rect -9473 747 -9439 781
rect -9281 747 -9247 781
rect -9089 747 -9055 781
rect -8897 747 -8863 781
rect -8705 747 -8671 781
rect -8513 747 -8479 781
rect -8321 747 -8287 781
rect -8129 747 -8095 781
rect -7937 747 -7903 781
rect -7745 747 -7711 781
rect -7553 747 -7519 781
rect -7361 747 -7327 781
rect -7169 747 -7135 781
rect -6977 747 -6943 781
rect -6785 747 -6751 781
rect -6593 747 -6559 781
rect -6401 747 -6367 781
rect -6209 747 -6175 781
rect -6017 747 -5983 781
rect -5825 747 -5791 781
rect -5633 747 -5599 781
rect -5441 747 -5407 781
rect -5249 747 -5215 781
rect -5057 747 -5023 781
rect -4865 747 -4831 781
rect -4673 747 -4639 781
rect -4481 747 -4447 781
rect -4289 747 -4255 781
rect -4097 747 -4063 781
rect -3905 747 -3871 781
rect -3713 747 -3679 781
rect -3521 747 -3487 781
rect -3329 747 -3295 781
rect -3137 747 -3103 781
rect -2945 747 -2911 781
rect -2753 747 -2719 781
rect -2561 747 -2527 781
rect -2369 747 -2335 781
rect -2177 747 -2143 781
rect -1985 747 -1951 781
rect -1793 747 -1759 781
rect -1601 747 -1567 781
rect -1409 747 -1375 781
rect -1217 747 -1183 781
rect -1025 747 -991 781
rect -833 747 -799 781
rect -641 747 -607 781
rect -449 747 -415 781
rect -257 747 -223 781
rect -65 747 -31 781
rect 127 747 161 781
rect 319 747 353 781
rect 511 747 545 781
rect 703 747 737 781
rect 895 747 929 781
rect 1087 747 1121 781
rect 1279 747 1313 781
rect 1471 747 1505 781
rect 1663 747 1697 781
rect 1855 747 1889 781
rect 2047 747 2081 781
rect 2239 747 2273 781
rect 2431 747 2465 781
rect 2623 747 2657 781
rect 2815 747 2849 781
rect 3007 747 3041 781
rect 3199 747 3233 781
rect 3391 747 3425 781
rect 3583 747 3617 781
rect 3775 747 3809 781
rect 3967 747 4001 781
rect 4159 747 4193 781
rect 4351 747 4385 781
rect 4543 747 4577 781
rect 4735 747 4769 781
rect 4927 747 4961 781
rect 5119 747 5153 781
rect 5311 747 5345 781
rect 5503 747 5537 781
rect 5695 747 5729 781
rect 5887 747 5921 781
rect 6079 747 6113 781
rect 6271 747 6305 781
rect 6463 747 6497 781
rect 6655 747 6689 781
rect 6847 747 6881 781
rect 7039 747 7073 781
rect 7231 747 7265 781
rect 7423 747 7457 781
rect 7615 747 7649 781
rect 7807 747 7841 781
rect 7999 747 8033 781
rect 8191 747 8225 781
rect 8383 747 8417 781
rect 8575 747 8609 781
rect 8767 747 8801 781
rect 8959 747 8993 781
rect 9151 747 9185 781
rect 9343 747 9377 781
rect 9535 747 9569 781
rect 9727 747 9761 781
rect 9919 747 9953 781
rect 10111 747 10145 781
rect 10303 747 10337 781
rect 10495 747 10529 781
rect -10577 -688 -10543 688
rect -10481 -688 -10447 688
rect -10385 -688 -10351 688
rect -10289 -688 -10255 688
rect -10193 -688 -10159 688
rect -10097 -688 -10063 688
rect -10001 -688 -9967 688
rect -9905 -688 -9871 688
rect -9809 -688 -9775 688
rect -9713 -688 -9679 688
rect -9617 -688 -9583 688
rect -9521 -688 -9487 688
rect -9425 -688 -9391 688
rect -9329 -688 -9295 688
rect -9233 -688 -9199 688
rect -9137 -688 -9103 688
rect -9041 -688 -9007 688
rect -8945 -688 -8911 688
rect -8849 -688 -8815 688
rect -8753 -688 -8719 688
rect -8657 -688 -8623 688
rect -8561 -688 -8527 688
rect -8465 -688 -8431 688
rect -8369 -688 -8335 688
rect -8273 -688 -8239 688
rect -8177 -688 -8143 688
rect -8081 -688 -8047 688
rect -7985 -688 -7951 688
rect -7889 -688 -7855 688
rect -7793 -688 -7759 688
rect -7697 -688 -7663 688
rect -7601 -688 -7567 688
rect -7505 -688 -7471 688
rect -7409 -688 -7375 688
rect -7313 -688 -7279 688
rect -7217 -688 -7183 688
rect -7121 -688 -7087 688
rect -7025 -688 -6991 688
rect -6929 -688 -6895 688
rect -6833 -688 -6799 688
rect -6737 -688 -6703 688
rect -6641 -688 -6607 688
rect -6545 -688 -6511 688
rect -6449 -688 -6415 688
rect -6353 -688 -6319 688
rect -6257 -688 -6223 688
rect -6161 -688 -6127 688
rect -6065 -688 -6031 688
rect -5969 -688 -5935 688
rect -5873 -688 -5839 688
rect -5777 -688 -5743 688
rect -5681 -688 -5647 688
rect -5585 -688 -5551 688
rect -5489 -688 -5455 688
rect -5393 -688 -5359 688
rect -5297 -688 -5263 688
rect -5201 -688 -5167 688
rect -5105 -688 -5071 688
rect -5009 -688 -4975 688
rect -4913 -688 -4879 688
rect -4817 -688 -4783 688
rect -4721 -688 -4687 688
rect -4625 -688 -4591 688
rect -4529 -688 -4495 688
rect -4433 -688 -4399 688
rect -4337 -688 -4303 688
rect -4241 -688 -4207 688
rect -4145 -688 -4111 688
rect -4049 -688 -4015 688
rect -3953 -688 -3919 688
rect -3857 -688 -3823 688
rect -3761 -688 -3727 688
rect -3665 -688 -3631 688
rect -3569 -688 -3535 688
rect -3473 -688 -3439 688
rect -3377 -688 -3343 688
rect -3281 -688 -3247 688
rect -3185 -688 -3151 688
rect -3089 -688 -3055 688
rect -2993 -688 -2959 688
rect -2897 -688 -2863 688
rect -2801 -688 -2767 688
rect -2705 -688 -2671 688
rect -2609 -688 -2575 688
rect -2513 -688 -2479 688
rect -2417 -688 -2383 688
rect -2321 -688 -2287 688
rect -2225 -688 -2191 688
rect -2129 -688 -2095 688
rect -2033 -688 -1999 688
rect -1937 -688 -1903 688
rect -1841 -688 -1807 688
rect -1745 -688 -1711 688
rect -1649 -688 -1615 688
rect -1553 -688 -1519 688
rect -1457 -688 -1423 688
rect -1361 -688 -1327 688
rect -1265 -688 -1231 688
rect -1169 -688 -1135 688
rect -1073 -688 -1039 688
rect -977 -688 -943 688
rect -881 -688 -847 688
rect -785 -688 -751 688
rect -689 -688 -655 688
rect -593 -688 -559 688
rect -497 -688 -463 688
rect -401 -688 -367 688
rect -305 -688 -271 688
rect -209 -688 -175 688
rect -113 -688 -79 688
rect -17 -688 17 688
rect 79 -688 113 688
rect 175 -688 209 688
rect 271 -688 305 688
rect 367 -688 401 688
rect 463 -688 497 688
rect 559 -688 593 688
rect 655 -688 689 688
rect 751 -688 785 688
rect 847 -688 881 688
rect 943 -688 977 688
rect 1039 -688 1073 688
rect 1135 -688 1169 688
rect 1231 -688 1265 688
rect 1327 -688 1361 688
rect 1423 -688 1457 688
rect 1519 -688 1553 688
rect 1615 -688 1649 688
rect 1711 -688 1745 688
rect 1807 -688 1841 688
rect 1903 -688 1937 688
rect 1999 -688 2033 688
rect 2095 -688 2129 688
rect 2191 -688 2225 688
rect 2287 -688 2321 688
rect 2383 -688 2417 688
rect 2479 -688 2513 688
rect 2575 -688 2609 688
rect 2671 -688 2705 688
rect 2767 -688 2801 688
rect 2863 -688 2897 688
rect 2959 -688 2993 688
rect 3055 -688 3089 688
rect 3151 -688 3185 688
rect 3247 -688 3281 688
rect 3343 -688 3377 688
rect 3439 -688 3473 688
rect 3535 -688 3569 688
rect 3631 -688 3665 688
rect 3727 -688 3761 688
rect 3823 -688 3857 688
rect 3919 -688 3953 688
rect 4015 -688 4049 688
rect 4111 -688 4145 688
rect 4207 -688 4241 688
rect 4303 -688 4337 688
rect 4399 -688 4433 688
rect 4495 -688 4529 688
rect 4591 -688 4625 688
rect 4687 -688 4721 688
rect 4783 -688 4817 688
rect 4879 -688 4913 688
rect 4975 -688 5009 688
rect 5071 -688 5105 688
rect 5167 -688 5201 688
rect 5263 -688 5297 688
rect 5359 -688 5393 688
rect 5455 -688 5489 688
rect 5551 -688 5585 688
rect 5647 -688 5681 688
rect 5743 -688 5777 688
rect 5839 -688 5873 688
rect 5935 -688 5969 688
rect 6031 -688 6065 688
rect 6127 -688 6161 688
rect 6223 -688 6257 688
rect 6319 -688 6353 688
rect 6415 -688 6449 688
rect 6511 -688 6545 688
rect 6607 -688 6641 688
rect 6703 -688 6737 688
rect 6799 -688 6833 688
rect 6895 -688 6929 688
rect 6991 -688 7025 688
rect 7087 -688 7121 688
rect 7183 -688 7217 688
rect 7279 -688 7313 688
rect 7375 -688 7409 688
rect 7471 -688 7505 688
rect 7567 -688 7601 688
rect 7663 -688 7697 688
rect 7759 -688 7793 688
rect 7855 -688 7889 688
rect 7951 -688 7985 688
rect 8047 -688 8081 688
rect 8143 -688 8177 688
rect 8239 -688 8273 688
rect 8335 -688 8369 688
rect 8431 -688 8465 688
rect 8527 -688 8561 688
rect 8623 -688 8657 688
rect 8719 -688 8753 688
rect 8815 -688 8849 688
rect 8911 -688 8945 688
rect 9007 -688 9041 688
rect 9103 -688 9137 688
rect 9199 -688 9233 688
rect 9295 -688 9329 688
rect 9391 -688 9425 688
rect 9487 -688 9521 688
rect 9583 -688 9617 688
rect 9679 -688 9713 688
rect 9775 -688 9809 688
rect 9871 -688 9905 688
rect 9967 -688 10001 688
rect 10063 -688 10097 688
rect 10159 -688 10193 688
rect 10255 -688 10289 688
rect 10351 -688 10385 688
rect 10447 -688 10481 688
rect 10543 -688 10577 688
rect -10529 -781 -10495 -747
rect -10337 -781 -10303 -747
rect -10145 -781 -10111 -747
rect -9953 -781 -9919 -747
rect -9761 -781 -9727 -747
rect -9569 -781 -9535 -747
rect -9377 -781 -9343 -747
rect -9185 -781 -9151 -747
rect -8993 -781 -8959 -747
rect -8801 -781 -8767 -747
rect -8609 -781 -8575 -747
rect -8417 -781 -8383 -747
rect -8225 -781 -8191 -747
rect -8033 -781 -7999 -747
rect -7841 -781 -7807 -747
rect -7649 -781 -7615 -747
rect -7457 -781 -7423 -747
rect -7265 -781 -7231 -747
rect -7073 -781 -7039 -747
rect -6881 -781 -6847 -747
rect -6689 -781 -6655 -747
rect -6497 -781 -6463 -747
rect -6305 -781 -6271 -747
rect -6113 -781 -6079 -747
rect -5921 -781 -5887 -747
rect -5729 -781 -5695 -747
rect -5537 -781 -5503 -747
rect -5345 -781 -5311 -747
rect -5153 -781 -5119 -747
rect -4961 -781 -4927 -747
rect -4769 -781 -4735 -747
rect -4577 -781 -4543 -747
rect -4385 -781 -4351 -747
rect -4193 -781 -4159 -747
rect -4001 -781 -3967 -747
rect -3809 -781 -3775 -747
rect -3617 -781 -3583 -747
rect -3425 -781 -3391 -747
rect -3233 -781 -3199 -747
rect -3041 -781 -3007 -747
rect -2849 -781 -2815 -747
rect -2657 -781 -2623 -747
rect -2465 -781 -2431 -747
rect -2273 -781 -2239 -747
rect -2081 -781 -2047 -747
rect -1889 -781 -1855 -747
rect -1697 -781 -1663 -747
rect -1505 -781 -1471 -747
rect -1313 -781 -1279 -747
rect -1121 -781 -1087 -747
rect -929 -781 -895 -747
rect -737 -781 -703 -747
rect -545 -781 -511 -747
rect -353 -781 -319 -747
rect -161 -781 -127 -747
rect 31 -781 65 -747
rect 223 -781 257 -747
rect 415 -781 449 -747
rect 607 -781 641 -747
rect 799 -781 833 -747
rect 991 -781 1025 -747
rect 1183 -781 1217 -747
rect 1375 -781 1409 -747
rect 1567 -781 1601 -747
rect 1759 -781 1793 -747
rect 1951 -781 1985 -747
rect 2143 -781 2177 -747
rect 2335 -781 2369 -747
rect 2527 -781 2561 -747
rect 2719 -781 2753 -747
rect 2911 -781 2945 -747
rect 3103 -781 3137 -747
rect 3295 -781 3329 -747
rect 3487 -781 3521 -747
rect 3679 -781 3713 -747
rect 3871 -781 3905 -747
rect 4063 -781 4097 -747
rect 4255 -781 4289 -747
rect 4447 -781 4481 -747
rect 4639 -781 4673 -747
rect 4831 -781 4865 -747
rect 5023 -781 5057 -747
rect 5215 -781 5249 -747
rect 5407 -781 5441 -747
rect 5599 -781 5633 -747
rect 5791 -781 5825 -747
rect 5983 -781 6017 -747
rect 6175 -781 6209 -747
rect 6367 -781 6401 -747
rect 6559 -781 6593 -747
rect 6751 -781 6785 -747
rect 6943 -781 6977 -747
rect 7135 -781 7169 -747
rect 7327 -781 7361 -747
rect 7519 -781 7553 -747
rect 7711 -781 7745 -747
rect 7903 -781 7937 -747
rect 8095 -781 8129 -747
rect 8287 -781 8321 -747
rect 8479 -781 8513 -747
rect 8671 -781 8705 -747
rect 8863 -781 8897 -747
rect 9055 -781 9089 -747
rect 9247 -781 9281 -747
rect 9439 -781 9473 -747
rect 9631 -781 9665 -747
rect 9823 -781 9857 -747
rect 10015 -781 10049 -747
rect 10207 -781 10241 -747
rect 10399 -781 10433 -747
<< metal1 >>
rect -10445 781 -10387 787
rect -10445 747 -10433 781
rect -10399 747 -10387 781
rect -10445 741 -10387 747
rect -10253 781 -10195 787
rect -10253 747 -10241 781
rect -10207 747 -10195 781
rect -10253 741 -10195 747
rect -10061 781 -10003 787
rect -10061 747 -10049 781
rect -10015 747 -10003 781
rect -10061 741 -10003 747
rect -9869 781 -9811 787
rect -9869 747 -9857 781
rect -9823 747 -9811 781
rect -9869 741 -9811 747
rect -9677 781 -9619 787
rect -9677 747 -9665 781
rect -9631 747 -9619 781
rect -9677 741 -9619 747
rect -9485 781 -9427 787
rect -9485 747 -9473 781
rect -9439 747 -9427 781
rect -9485 741 -9427 747
rect -9293 781 -9235 787
rect -9293 747 -9281 781
rect -9247 747 -9235 781
rect -9293 741 -9235 747
rect -9101 781 -9043 787
rect -9101 747 -9089 781
rect -9055 747 -9043 781
rect -9101 741 -9043 747
rect -8909 781 -8851 787
rect -8909 747 -8897 781
rect -8863 747 -8851 781
rect -8909 741 -8851 747
rect -8717 781 -8659 787
rect -8717 747 -8705 781
rect -8671 747 -8659 781
rect -8717 741 -8659 747
rect -8525 781 -8467 787
rect -8525 747 -8513 781
rect -8479 747 -8467 781
rect -8525 741 -8467 747
rect -8333 781 -8275 787
rect -8333 747 -8321 781
rect -8287 747 -8275 781
rect -8333 741 -8275 747
rect -8141 781 -8083 787
rect -8141 747 -8129 781
rect -8095 747 -8083 781
rect -8141 741 -8083 747
rect -7949 781 -7891 787
rect -7949 747 -7937 781
rect -7903 747 -7891 781
rect -7949 741 -7891 747
rect -7757 781 -7699 787
rect -7757 747 -7745 781
rect -7711 747 -7699 781
rect -7757 741 -7699 747
rect -7565 781 -7507 787
rect -7565 747 -7553 781
rect -7519 747 -7507 781
rect -7565 741 -7507 747
rect -7373 781 -7315 787
rect -7373 747 -7361 781
rect -7327 747 -7315 781
rect -7373 741 -7315 747
rect -7181 781 -7123 787
rect -7181 747 -7169 781
rect -7135 747 -7123 781
rect -7181 741 -7123 747
rect -6989 781 -6931 787
rect -6989 747 -6977 781
rect -6943 747 -6931 781
rect -6989 741 -6931 747
rect -6797 781 -6739 787
rect -6797 747 -6785 781
rect -6751 747 -6739 781
rect -6797 741 -6739 747
rect -6605 781 -6547 787
rect -6605 747 -6593 781
rect -6559 747 -6547 781
rect -6605 741 -6547 747
rect -6413 781 -6355 787
rect -6413 747 -6401 781
rect -6367 747 -6355 781
rect -6413 741 -6355 747
rect -6221 781 -6163 787
rect -6221 747 -6209 781
rect -6175 747 -6163 781
rect -6221 741 -6163 747
rect -6029 781 -5971 787
rect -6029 747 -6017 781
rect -5983 747 -5971 781
rect -6029 741 -5971 747
rect -5837 781 -5779 787
rect -5837 747 -5825 781
rect -5791 747 -5779 781
rect -5837 741 -5779 747
rect -5645 781 -5587 787
rect -5645 747 -5633 781
rect -5599 747 -5587 781
rect -5645 741 -5587 747
rect -5453 781 -5395 787
rect -5453 747 -5441 781
rect -5407 747 -5395 781
rect -5453 741 -5395 747
rect -5261 781 -5203 787
rect -5261 747 -5249 781
rect -5215 747 -5203 781
rect -5261 741 -5203 747
rect -5069 781 -5011 787
rect -5069 747 -5057 781
rect -5023 747 -5011 781
rect -5069 741 -5011 747
rect -4877 781 -4819 787
rect -4877 747 -4865 781
rect -4831 747 -4819 781
rect -4877 741 -4819 747
rect -4685 781 -4627 787
rect -4685 747 -4673 781
rect -4639 747 -4627 781
rect -4685 741 -4627 747
rect -4493 781 -4435 787
rect -4493 747 -4481 781
rect -4447 747 -4435 781
rect -4493 741 -4435 747
rect -4301 781 -4243 787
rect -4301 747 -4289 781
rect -4255 747 -4243 781
rect -4301 741 -4243 747
rect -4109 781 -4051 787
rect -4109 747 -4097 781
rect -4063 747 -4051 781
rect -4109 741 -4051 747
rect -3917 781 -3859 787
rect -3917 747 -3905 781
rect -3871 747 -3859 781
rect -3917 741 -3859 747
rect -3725 781 -3667 787
rect -3725 747 -3713 781
rect -3679 747 -3667 781
rect -3725 741 -3667 747
rect -3533 781 -3475 787
rect -3533 747 -3521 781
rect -3487 747 -3475 781
rect -3533 741 -3475 747
rect -3341 781 -3283 787
rect -3341 747 -3329 781
rect -3295 747 -3283 781
rect -3341 741 -3283 747
rect -3149 781 -3091 787
rect -3149 747 -3137 781
rect -3103 747 -3091 781
rect -3149 741 -3091 747
rect -2957 781 -2899 787
rect -2957 747 -2945 781
rect -2911 747 -2899 781
rect -2957 741 -2899 747
rect -2765 781 -2707 787
rect -2765 747 -2753 781
rect -2719 747 -2707 781
rect -2765 741 -2707 747
rect -2573 781 -2515 787
rect -2573 747 -2561 781
rect -2527 747 -2515 781
rect -2573 741 -2515 747
rect -2381 781 -2323 787
rect -2381 747 -2369 781
rect -2335 747 -2323 781
rect -2381 741 -2323 747
rect -2189 781 -2131 787
rect -2189 747 -2177 781
rect -2143 747 -2131 781
rect -2189 741 -2131 747
rect -1997 781 -1939 787
rect -1997 747 -1985 781
rect -1951 747 -1939 781
rect -1997 741 -1939 747
rect -1805 781 -1747 787
rect -1805 747 -1793 781
rect -1759 747 -1747 781
rect -1805 741 -1747 747
rect -1613 781 -1555 787
rect -1613 747 -1601 781
rect -1567 747 -1555 781
rect -1613 741 -1555 747
rect -1421 781 -1363 787
rect -1421 747 -1409 781
rect -1375 747 -1363 781
rect -1421 741 -1363 747
rect -1229 781 -1171 787
rect -1229 747 -1217 781
rect -1183 747 -1171 781
rect -1229 741 -1171 747
rect -1037 781 -979 787
rect -1037 747 -1025 781
rect -991 747 -979 781
rect -1037 741 -979 747
rect -845 781 -787 787
rect -845 747 -833 781
rect -799 747 -787 781
rect -845 741 -787 747
rect -653 781 -595 787
rect -653 747 -641 781
rect -607 747 -595 781
rect -653 741 -595 747
rect -461 781 -403 787
rect -461 747 -449 781
rect -415 747 -403 781
rect -461 741 -403 747
rect -269 781 -211 787
rect -269 747 -257 781
rect -223 747 -211 781
rect -269 741 -211 747
rect -77 781 -19 787
rect -77 747 -65 781
rect -31 747 -19 781
rect -77 741 -19 747
rect 115 781 173 787
rect 115 747 127 781
rect 161 747 173 781
rect 115 741 173 747
rect 307 781 365 787
rect 307 747 319 781
rect 353 747 365 781
rect 307 741 365 747
rect 499 781 557 787
rect 499 747 511 781
rect 545 747 557 781
rect 499 741 557 747
rect 691 781 749 787
rect 691 747 703 781
rect 737 747 749 781
rect 691 741 749 747
rect 883 781 941 787
rect 883 747 895 781
rect 929 747 941 781
rect 883 741 941 747
rect 1075 781 1133 787
rect 1075 747 1087 781
rect 1121 747 1133 781
rect 1075 741 1133 747
rect 1267 781 1325 787
rect 1267 747 1279 781
rect 1313 747 1325 781
rect 1267 741 1325 747
rect 1459 781 1517 787
rect 1459 747 1471 781
rect 1505 747 1517 781
rect 1459 741 1517 747
rect 1651 781 1709 787
rect 1651 747 1663 781
rect 1697 747 1709 781
rect 1651 741 1709 747
rect 1843 781 1901 787
rect 1843 747 1855 781
rect 1889 747 1901 781
rect 1843 741 1901 747
rect 2035 781 2093 787
rect 2035 747 2047 781
rect 2081 747 2093 781
rect 2035 741 2093 747
rect 2227 781 2285 787
rect 2227 747 2239 781
rect 2273 747 2285 781
rect 2227 741 2285 747
rect 2419 781 2477 787
rect 2419 747 2431 781
rect 2465 747 2477 781
rect 2419 741 2477 747
rect 2611 781 2669 787
rect 2611 747 2623 781
rect 2657 747 2669 781
rect 2611 741 2669 747
rect 2803 781 2861 787
rect 2803 747 2815 781
rect 2849 747 2861 781
rect 2803 741 2861 747
rect 2995 781 3053 787
rect 2995 747 3007 781
rect 3041 747 3053 781
rect 2995 741 3053 747
rect 3187 781 3245 787
rect 3187 747 3199 781
rect 3233 747 3245 781
rect 3187 741 3245 747
rect 3379 781 3437 787
rect 3379 747 3391 781
rect 3425 747 3437 781
rect 3379 741 3437 747
rect 3571 781 3629 787
rect 3571 747 3583 781
rect 3617 747 3629 781
rect 3571 741 3629 747
rect 3763 781 3821 787
rect 3763 747 3775 781
rect 3809 747 3821 781
rect 3763 741 3821 747
rect 3955 781 4013 787
rect 3955 747 3967 781
rect 4001 747 4013 781
rect 3955 741 4013 747
rect 4147 781 4205 787
rect 4147 747 4159 781
rect 4193 747 4205 781
rect 4147 741 4205 747
rect 4339 781 4397 787
rect 4339 747 4351 781
rect 4385 747 4397 781
rect 4339 741 4397 747
rect 4531 781 4589 787
rect 4531 747 4543 781
rect 4577 747 4589 781
rect 4531 741 4589 747
rect 4723 781 4781 787
rect 4723 747 4735 781
rect 4769 747 4781 781
rect 4723 741 4781 747
rect 4915 781 4973 787
rect 4915 747 4927 781
rect 4961 747 4973 781
rect 4915 741 4973 747
rect 5107 781 5165 787
rect 5107 747 5119 781
rect 5153 747 5165 781
rect 5107 741 5165 747
rect 5299 781 5357 787
rect 5299 747 5311 781
rect 5345 747 5357 781
rect 5299 741 5357 747
rect 5491 781 5549 787
rect 5491 747 5503 781
rect 5537 747 5549 781
rect 5491 741 5549 747
rect 5683 781 5741 787
rect 5683 747 5695 781
rect 5729 747 5741 781
rect 5683 741 5741 747
rect 5875 781 5933 787
rect 5875 747 5887 781
rect 5921 747 5933 781
rect 5875 741 5933 747
rect 6067 781 6125 787
rect 6067 747 6079 781
rect 6113 747 6125 781
rect 6067 741 6125 747
rect 6259 781 6317 787
rect 6259 747 6271 781
rect 6305 747 6317 781
rect 6259 741 6317 747
rect 6451 781 6509 787
rect 6451 747 6463 781
rect 6497 747 6509 781
rect 6451 741 6509 747
rect 6643 781 6701 787
rect 6643 747 6655 781
rect 6689 747 6701 781
rect 6643 741 6701 747
rect 6835 781 6893 787
rect 6835 747 6847 781
rect 6881 747 6893 781
rect 6835 741 6893 747
rect 7027 781 7085 787
rect 7027 747 7039 781
rect 7073 747 7085 781
rect 7027 741 7085 747
rect 7219 781 7277 787
rect 7219 747 7231 781
rect 7265 747 7277 781
rect 7219 741 7277 747
rect 7411 781 7469 787
rect 7411 747 7423 781
rect 7457 747 7469 781
rect 7411 741 7469 747
rect 7603 781 7661 787
rect 7603 747 7615 781
rect 7649 747 7661 781
rect 7603 741 7661 747
rect 7795 781 7853 787
rect 7795 747 7807 781
rect 7841 747 7853 781
rect 7795 741 7853 747
rect 7987 781 8045 787
rect 7987 747 7999 781
rect 8033 747 8045 781
rect 7987 741 8045 747
rect 8179 781 8237 787
rect 8179 747 8191 781
rect 8225 747 8237 781
rect 8179 741 8237 747
rect 8371 781 8429 787
rect 8371 747 8383 781
rect 8417 747 8429 781
rect 8371 741 8429 747
rect 8563 781 8621 787
rect 8563 747 8575 781
rect 8609 747 8621 781
rect 8563 741 8621 747
rect 8755 781 8813 787
rect 8755 747 8767 781
rect 8801 747 8813 781
rect 8755 741 8813 747
rect 8947 781 9005 787
rect 8947 747 8959 781
rect 8993 747 9005 781
rect 8947 741 9005 747
rect 9139 781 9197 787
rect 9139 747 9151 781
rect 9185 747 9197 781
rect 9139 741 9197 747
rect 9331 781 9389 787
rect 9331 747 9343 781
rect 9377 747 9389 781
rect 9331 741 9389 747
rect 9523 781 9581 787
rect 9523 747 9535 781
rect 9569 747 9581 781
rect 9523 741 9581 747
rect 9715 781 9773 787
rect 9715 747 9727 781
rect 9761 747 9773 781
rect 9715 741 9773 747
rect 9907 781 9965 787
rect 9907 747 9919 781
rect 9953 747 9965 781
rect 9907 741 9965 747
rect 10099 781 10157 787
rect 10099 747 10111 781
rect 10145 747 10157 781
rect 10099 741 10157 747
rect 10291 781 10349 787
rect 10291 747 10303 781
rect 10337 747 10349 781
rect 10291 741 10349 747
rect 10483 781 10541 787
rect 10483 747 10495 781
rect 10529 747 10541 781
rect 10483 741 10541 747
rect -10583 688 -10537 700
rect -10583 -688 -10577 688
rect -10543 -688 -10537 688
rect -10583 -700 -10537 -688
rect -10487 688 -10441 700
rect -10487 -688 -10481 688
rect -10447 -688 -10441 688
rect -10487 -700 -10441 -688
rect -10391 688 -10345 700
rect -10391 -688 -10385 688
rect -10351 -688 -10345 688
rect -10391 -700 -10345 -688
rect -10295 688 -10249 700
rect -10295 -688 -10289 688
rect -10255 -688 -10249 688
rect -10295 -700 -10249 -688
rect -10199 688 -10153 700
rect -10199 -688 -10193 688
rect -10159 -688 -10153 688
rect -10199 -700 -10153 -688
rect -10103 688 -10057 700
rect -10103 -688 -10097 688
rect -10063 -688 -10057 688
rect -10103 -700 -10057 -688
rect -10007 688 -9961 700
rect -10007 -688 -10001 688
rect -9967 -688 -9961 688
rect -10007 -700 -9961 -688
rect -9911 688 -9865 700
rect -9911 -688 -9905 688
rect -9871 -688 -9865 688
rect -9911 -700 -9865 -688
rect -9815 688 -9769 700
rect -9815 -688 -9809 688
rect -9775 -688 -9769 688
rect -9815 -700 -9769 -688
rect -9719 688 -9673 700
rect -9719 -688 -9713 688
rect -9679 -688 -9673 688
rect -9719 -700 -9673 -688
rect -9623 688 -9577 700
rect -9623 -688 -9617 688
rect -9583 -688 -9577 688
rect -9623 -700 -9577 -688
rect -9527 688 -9481 700
rect -9527 -688 -9521 688
rect -9487 -688 -9481 688
rect -9527 -700 -9481 -688
rect -9431 688 -9385 700
rect -9431 -688 -9425 688
rect -9391 -688 -9385 688
rect -9431 -700 -9385 -688
rect -9335 688 -9289 700
rect -9335 -688 -9329 688
rect -9295 -688 -9289 688
rect -9335 -700 -9289 -688
rect -9239 688 -9193 700
rect -9239 -688 -9233 688
rect -9199 -688 -9193 688
rect -9239 -700 -9193 -688
rect -9143 688 -9097 700
rect -9143 -688 -9137 688
rect -9103 -688 -9097 688
rect -9143 -700 -9097 -688
rect -9047 688 -9001 700
rect -9047 -688 -9041 688
rect -9007 -688 -9001 688
rect -9047 -700 -9001 -688
rect -8951 688 -8905 700
rect -8951 -688 -8945 688
rect -8911 -688 -8905 688
rect -8951 -700 -8905 -688
rect -8855 688 -8809 700
rect -8855 -688 -8849 688
rect -8815 -688 -8809 688
rect -8855 -700 -8809 -688
rect -8759 688 -8713 700
rect -8759 -688 -8753 688
rect -8719 -688 -8713 688
rect -8759 -700 -8713 -688
rect -8663 688 -8617 700
rect -8663 -688 -8657 688
rect -8623 -688 -8617 688
rect -8663 -700 -8617 -688
rect -8567 688 -8521 700
rect -8567 -688 -8561 688
rect -8527 -688 -8521 688
rect -8567 -700 -8521 -688
rect -8471 688 -8425 700
rect -8471 -688 -8465 688
rect -8431 -688 -8425 688
rect -8471 -700 -8425 -688
rect -8375 688 -8329 700
rect -8375 -688 -8369 688
rect -8335 -688 -8329 688
rect -8375 -700 -8329 -688
rect -8279 688 -8233 700
rect -8279 -688 -8273 688
rect -8239 -688 -8233 688
rect -8279 -700 -8233 -688
rect -8183 688 -8137 700
rect -8183 -688 -8177 688
rect -8143 -688 -8137 688
rect -8183 -700 -8137 -688
rect -8087 688 -8041 700
rect -8087 -688 -8081 688
rect -8047 -688 -8041 688
rect -8087 -700 -8041 -688
rect -7991 688 -7945 700
rect -7991 -688 -7985 688
rect -7951 -688 -7945 688
rect -7991 -700 -7945 -688
rect -7895 688 -7849 700
rect -7895 -688 -7889 688
rect -7855 -688 -7849 688
rect -7895 -700 -7849 -688
rect -7799 688 -7753 700
rect -7799 -688 -7793 688
rect -7759 -688 -7753 688
rect -7799 -700 -7753 -688
rect -7703 688 -7657 700
rect -7703 -688 -7697 688
rect -7663 -688 -7657 688
rect -7703 -700 -7657 -688
rect -7607 688 -7561 700
rect -7607 -688 -7601 688
rect -7567 -688 -7561 688
rect -7607 -700 -7561 -688
rect -7511 688 -7465 700
rect -7511 -688 -7505 688
rect -7471 -688 -7465 688
rect -7511 -700 -7465 -688
rect -7415 688 -7369 700
rect -7415 -688 -7409 688
rect -7375 -688 -7369 688
rect -7415 -700 -7369 -688
rect -7319 688 -7273 700
rect -7319 -688 -7313 688
rect -7279 -688 -7273 688
rect -7319 -700 -7273 -688
rect -7223 688 -7177 700
rect -7223 -688 -7217 688
rect -7183 -688 -7177 688
rect -7223 -700 -7177 -688
rect -7127 688 -7081 700
rect -7127 -688 -7121 688
rect -7087 -688 -7081 688
rect -7127 -700 -7081 -688
rect -7031 688 -6985 700
rect -7031 -688 -7025 688
rect -6991 -688 -6985 688
rect -7031 -700 -6985 -688
rect -6935 688 -6889 700
rect -6935 -688 -6929 688
rect -6895 -688 -6889 688
rect -6935 -700 -6889 -688
rect -6839 688 -6793 700
rect -6839 -688 -6833 688
rect -6799 -688 -6793 688
rect -6839 -700 -6793 -688
rect -6743 688 -6697 700
rect -6743 -688 -6737 688
rect -6703 -688 -6697 688
rect -6743 -700 -6697 -688
rect -6647 688 -6601 700
rect -6647 -688 -6641 688
rect -6607 -688 -6601 688
rect -6647 -700 -6601 -688
rect -6551 688 -6505 700
rect -6551 -688 -6545 688
rect -6511 -688 -6505 688
rect -6551 -700 -6505 -688
rect -6455 688 -6409 700
rect -6455 -688 -6449 688
rect -6415 -688 -6409 688
rect -6455 -700 -6409 -688
rect -6359 688 -6313 700
rect -6359 -688 -6353 688
rect -6319 -688 -6313 688
rect -6359 -700 -6313 -688
rect -6263 688 -6217 700
rect -6263 -688 -6257 688
rect -6223 -688 -6217 688
rect -6263 -700 -6217 -688
rect -6167 688 -6121 700
rect -6167 -688 -6161 688
rect -6127 -688 -6121 688
rect -6167 -700 -6121 -688
rect -6071 688 -6025 700
rect -6071 -688 -6065 688
rect -6031 -688 -6025 688
rect -6071 -700 -6025 -688
rect -5975 688 -5929 700
rect -5975 -688 -5969 688
rect -5935 -688 -5929 688
rect -5975 -700 -5929 -688
rect -5879 688 -5833 700
rect -5879 -688 -5873 688
rect -5839 -688 -5833 688
rect -5879 -700 -5833 -688
rect -5783 688 -5737 700
rect -5783 -688 -5777 688
rect -5743 -688 -5737 688
rect -5783 -700 -5737 -688
rect -5687 688 -5641 700
rect -5687 -688 -5681 688
rect -5647 -688 -5641 688
rect -5687 -700 -5641 -688
rect -5591 688 -5545 700
rect -5591 -688 -5585 688
rect -5551 -688 -5545 688
rect -5591 -700 -5545 -688
rect -5495 688 -5449 700
rect -5495 -688 -5489 688
rect -5455 -688 -5449 688
rect -5495 -700 -5449 -688
rect -5399 688 -5353 700
rect -5399 -688 -5393 688
rect -5359 -688 -5353 688
rect -5399 -700 -5353 -688
rect -5303 688 -5257 700
rect -5303 -688 -5297 688
rect -5263 -688 -5257 688
rect -5303 -700 -5257 -688
rect -5207 688 -5161 700
rect -5207 -688 -5201 688
rect -5167 -688 -5161 688
rect -5207 -700 -5161 -688
rect -5111 688 -5065 700
rect -5111 -688 -5105 688
rect -5071 -688 -5065 688
rect -5111 -700 -5065 -688
rect -5015 688 -4969 700
rect -5015 -688 -5009 688
rect -4975 -688 -4969 688
rect -5015 -700 -4969 -688
rect -4919 688 -4873 700
rect -4919 -688 -4913 688
rect -4879 -688 -4873 688
rect -4919 -700 -4873 -688
rect -4823 688 -4777 700
rect -4823 -688 -4817 688
rect -4783 -688 -4777 688
rect -4823 -700 -4777 -688
rect -4727 688 -4681 700
rect -4727 -688 -4721 688
rect -4687 -688 -4681 688
rect -4727 -700 -4681 -688
rect -4631 688 -4585 700
rect -4631 -688 -4625 688
rect -4591 -688 -4585 688
rect -4631 -700 -4585 -688
rect -4535 688 -4489 700
rect -4535 -688 -4529 688
rect -4495 -688 -4489 688
rect -4535 -700 -4489 -688
rect -4439 688 -4393 700
rect -4439 -688 -4433 688
rect -4399 -688 -4393 688
rect -4439 -700 -4393 -688
rect -4343 688 -4297 700
rect -4343 -688 -4337 688
rect -4303 -688 -4297 688
rect -4343 -700 -4297 -688
rect -4247 688 -4201 700
rect -4247 -688 -4241 688
rect -4207 -688 -4201 688
rect -4247 -700 -4201 -688
rect -4151 688 -4105 700
rect -4151 -688 -4145 688
rect -4111 -688 -4105 688
rect -4151 -700 -4105 -688
rect -4055 688 -4009 700
rect -4055 -688 -4049 688
rect -4015 -688 -4009 688
rect -4055 -700 -4009 -688
rect -3959 688 -3913 700
rect -3959 -688 -3953 688
rect -3919 -688 -3913 688
rect -3959 -700 -3913 -688
rect -3863 688 -3817 700
rect -3863 -688 -3857 688
rect -3823 -688 -3817 688
rect -3863 -700 -3817 -688
rect -3767 688 -3721 700
rect -3767 -688 -3761 688
rect -3727 -688 -3721 688
rect -3767 -700 -3721 -688
rect -3671 688 -3625 700
rect -3671 -688 -3665 688
rect -3631 -688 -3625 688
rect -3671 -700 -3625 -688
rect -3575 688 -3529 700
rect -3575 -688 -3569 688
rect -3535 -688 -3529 688
rect -3575 -700 -3529 -688
rect -3479 688 -3433 700
rect -3479 -688 -3473 688
rect -3439 -688 -3433 688
rect -3479 -700 -3433 -688
rect -3383 688 -3337 700
rect -3383 -688 -3377 688
rect -3343 -688 -3337 688
rect -3383 -700 -3337 -688
rect -3287 688 -3241 700
rect -3287 -688 -3281 688
rect -3247 -688 -3241 688
rect -3287 -700 -3241 -688
rect -3191 688 -3145 700
rect -3191 -688 -3185 688
rect -3151 -688 -3145 688
rect -3191 -700 -3145 -688
rect -3095 688 -3049 700
rect -3095 -688 -3089 688
rect -3055 -688 -3049 688
rect -3095 -700 -3049 -688
rect -2999 688 -2953 700
rect -2999 -688 -2993 688
rect -2959 -688 -2953 688
rect -2999 -700 -2953 -688
rect -2903 688 -2857 700
rect -2903 -688 -2897 688
rect -2863 -688 -2857 688
rect -2903 -700 -2857 -688
rect -2807 688 -2761 700
rect -2807 -688 -2801 688
rect -2767 -688 -2761 688
rect -2807 -700 -2761 -688
rect -2711 688 -2665 700
rect -2711 -688 -2705 688
rect -2671 -688 -2665 688
rect -2711 -700 -2665 -688
rect -2615 688 -2569 700
rect -2615 -688 -2609 688
rect -2575 -688 -2569 688
rect -2615 -700 -2569 -688
rect -2519 688 -2473 700
rect -2519 -688 -2513 688
rect -2479 -688 -2473 688
rect -2519 -700 -2473 -688
rect -2423 688 -2377 700
rect -2423 -688 -2417 688
rect -2383 -688 -2377 688
rect -2423 -700 -2377 -688
rect -2327 688 -2281 700
rect -2327 -688 -2321 688
rect -2287 -688 -2281 688
rect -2327 -700 -2281 -688
rect -2231 688 -2185 700
rect -2231 -688 -2225 688
rect -2191 -688 -2185 688
rect -2231 -700 -2185 -688
rect -2135 688 -2089 700
rect -2135 -688 -2129 688
rect -2095 -688 -2089 688
rect -2135 -700 -2089 -688
rect -2039 688 -1993 700
rect -2039 -688 -2033 688
rect -1999 -688 -1993 688
rect -2039 -700 -1993 -688
rect -1943 688 -1897 700
rect -1943 -688 -1937 688
rect -1903 -688 -1897 688
rect -1943 -700 -1897 -688
rect -1847 688 -1801 700
rect -1847 -688 -1841 688
rect -1807 -688 -1801 688
rect -1847 -700 -1801 -688
rect -1751 688 -1705 700
rect -1751 -688 -1745 688
rect -1711 -688 -1705 688
rect -1751 -700 -1705 -688
rect -1655 688 -1609 700
rect -1655 -688 -1649 688
rect -1615 -688 -1609 688
rect -1655 -700 -1609 -688
rect -1559 688 -1513 700
rect -1559 -688 -1553 688
rect -1519 -688 -1513 688
rect -1559 -700 -1513 -688
rect -1463 688 -1417 700
rect -1463 -688 -1457 688
rect -1423 -688 -1417 688
rect -1463 -700 -1417 -688
rect -1367 688 -1321 700
rect -1367 -688 -1361 688
rect -1327 -688 -1321 688
rect -1367 -700 -1321 -688
rect -1271 688 -1225 700
rect -1271 -688 -1265 688
rect -1231 -688 -1225 688
rect -1271 -700 -1225 -688
rect -1175 688 -1129 700
rect -1175 -688 -1169 688
rect -1135 -688 -1129 688
rect -1175 -700 -1129 -688
rect -1079 688 -1033 700
rect -1079 -688 -1073 688
rect -1039 -688 -1033 688
rect -1079 -700 -1033 -688
rect -983 688 -937 700
rect -983 -688 -977 688
rect -943 -688 -937 688
rect -983 -700 -937 -688
rect -887 688 -841 700
rect -887 -688 -881 688
rect -847 -688 -841 688
rect -887 -700 -841 -688
rect -791 688 -745 700
rect -791 -688 -785 688
rect -751 -688 -745 688
rect -791 -700 -745 -688
rect -695 688 -649 700
rect -695 -688 -689 688
rect -655 -688 -649 688
rect -695 -700 -649 -688
rect -599 688 -553 700
rect -599 -688 -593 688
rect -559 -688 -553 688
rect -599 -700 -553 -688
rect -503 688 -457 700
rect -503 -688 -497 688
rect -463 -688 -457 688
rect -503 -700 -457 -688
rect -407 688 -361 700
rect -407 -688 -401 688
rect -367 -688 -361 688
rect -407 -700 -361 -688
rect -311 688 -265 700
rect -311 -688 -305 688
rect -271 -688 -265 688
rect -311 -700 -265 -688
rect -215 688 -169 700
rect -215 -688 -209 688
rect -175 -688 -169 688
rect -215 -700 -169 -688
rect -119 688 -73 700
rect -119 -688 -113 688
rect -79 -688 -73 688
rect -119 -700 -73 -688
rect -23 688 23 700
rect -23 -688 -17 688
rect 17 -688 23 688
rect -23 -700 23 -688
rect 73 688 119 700
rect 73 -688 79 688
rect 113 -688 119 688
rect 73 -700 119 -688
rect 169 688 215 700
rect 169 -688 175 688
rect 209 -688 215 688
rect 169 -700 215 -688
rect 265 688 311 700
rect 265 -688 271 688
rect 305 -688 311 688
rect 265 -700 311 -688
rect 361 688 407 700
rect 361 -688 367 688
rect 401 -688 407 688
rect 361 -700 407 -688
rect 457 688 503 700
rect 457 -688 463 688
rect 497 -688 503 688
rect 457 -700 503 -688
rect 553 688 599 700
rect 553 -688 559 688
rect 593 -688 599 688
rect 553 -700 599 -688
rect 649 688 695 700
rect 649 -688 655 688
rect 689 -688 695 688
rect 649 -700 695 -688
rect 745 688 791 700
rect 745 -688 751 688
rect 785 -688 791 688
rect 745 -700 791 -688
rect 841 688 887 700
rect 841 -688 847 688
rect 881 -688 887 688
rect 841 -700 887 -688
rect 937 688 983 700
rect 937 -688 943 688
rect 977 -688 983 688
rect 937 -700 983 -688
rect 1033 688 1079 700
rect 1033 -688 1039 688
rect 1073 -688 1079 688
rect 1033 -700 1079 -688
rect 1129 688 1175 700
rect 1129 -688 1135 688
rect 1169 -688 1175 688
rect 1129 -700 1175 -688
rect 1225 688 1271 700
rect 1225 -688 1231 688
rect 1265 -688 1271 688
rect 1225 -700 1271 -688
rect 1321 688 1367 700
rect 1321 -688 1327 688
rect 1361 -688 1367 688
rect 1321 -700 1367 -688
rect 1417 688 1463 700
rect 1417 -688 1423 688
rect 1457 -688 1463 688
rect 1417 -700 1463 -688
rect 1513 688 1559 700
rect 1513 -688 1519 688
rect 1553 -688 1559 688
rect 1513 -700 1559 -688
rect 1609 688 1655 700
rect 1609 -688 1615 688
rect 1649 -688 1655 688
rect 1609 -700 1655 -688
rect 1705 688 1751 700
rect 1705 -688 1711 688
rect 1745 -688 1751 688
rect 1705 -700 1751 -688
rect 1801 688 1847 700
rect 1801 -688 1807 688
rect 1841 -688 1847 688
rect 1801 -700 1847 -688
rect 1897 688 1943 700
rect 1897 -688 1903 688
rect 1937 -688 1943 688
rect 1897 -700 1943 -688
rect 1993 688 2039 700
rect 1993 -688 1999 688
rect 2033 -688 2039 688
rect 1993 -700 2039 -688
rect 2089 688 2135 700
rect 2089 -688 2095 688
rect 2129 -688 2135 688
rect 2089 -700 2135 -688
rect 2185 688 2231 700
rect 2185 -688 2191 688
rect 2225 -688 2231 688
rect 2185 -700 2231 -688
rect 2281 688 2327 700
rect 2281 -688 2287 688
rect 2321 -688 2327 688
rect 2281 -700 2327 -688
rect 2377 688 2423 700
rect 2377 -688 2383 688
rect 2417 -688 2423 688
rect 2377 -700 2423 -688
rect 2473 688 2519 700
rect 2473 -688 2479 688
rect 2513 -688 2519 688
rect 2473 -700 2519 -688
rect 2569 688 2615 700
rect 2569 -688 2575 688
rect 2609 -688 2615 688
rect 2569 -700 2615 -688
rect 2665 688 2711 700
rect 2665 -688 2671 688
rect 2705 -688 2711 688
rect 2665 -700 2711 -688
rect 2761 688 2807 700
rect 2761 -688 2767 688
rect 2801 -688 2807 688
rect 2761 -700 2807 -688
rect 2857 688 2903 700
rect 2857 -688 2863 688
rect 2897 -688 2903 688
rect 2857 -700 2903 -688
rect 2953 688 2999 700
rect 2953 -688 2959 688
rect 2993 -688 2999 688
rect 2953 -700 2999 -688
rect 3049 688 3095 700
rect 3049 -688 3055 688
rect 3089 -688 3095 688
rect 3049 -700 3095 -688
rect 3145 688 3191 700
rect 3145 -688 3151 688
rect 3185 -688 3191 688
rect 3145 -700 3191 -688
rect 3241 688 3287 700
rect 3241 -688 3247 688
rect 3281 -688 3287 688
rect 3241 -700 3287 -688
rect 3337 688 3383 700
rect 3337 -688 3343 688
rect 3377 -688 3383 688
rect 3337 -700 3383 -688
rect 3433 688 3479 700
rect 3433 -688 3439 688
rect 3473 -688 3479 688
rect 3433 -700 3479 -688
rect 3529 688 3575 700
rect 3529 -688 3535 688
rect 3569 -688 3575 688
rect 3529 -700 3575 -688
rect 3625 688 3671 700
rect 3625 -688 3631 688
rect 3665 -688 3671 688
rect 3625 -700 3671 -688
rect 3721 688 3767 700
rect 3721 -688 3727 688
rect 3761 -688 3767 688
rect 3721 -700 3767 -688
rect 3817 688 3863 700
rect 3817 -688 3823 688
rect 3857 -688 3863 688
rect 3817 -700 3863 -688
rect 3913 688 3959 700
rect 3913 -688 3919 688
rect 3953 -688 3959 688
rect 3913 -700 3959 -688
rect 4009 688 4055 700
rect 4009 -688 4015 688
rect 4049 -688 4055 688
rect 4009 -700 4055 -688
rect 4105 688 4151 700
rect 4105 -688 4111 688
rect 4145 -688 4151 688
rect 4105 -700 4151 -688
rect 4201 688 4247 700
rect 4201 -688 4207 688
rect 4241 -688 4247 688
rect 4201 -700 4247 -688
rect 4297 688 4343 700
rect 4297 -688 4303 688
rect 4337 -688 4343 688
rect 4297 -700 4343 -688
rect 4393 688 4439 700
rect 4393 -688 4399 688
rect 4433 -688 4439 688
rect 4393 -700 4439 -688
rect 4489 688 4535 700
rect 4489 -688 4495 688
rect 4529 -688 4535 688
rect 4489 -700 4535 -688
rect 4585 688 4631 700
rect 4585 -688 4591 688
rect 4625 -688 4631 688
rect 4585 -700 4631 -688
rect 4681 688 4727 700
rect 4681 -688 4687 688
rect 4721 -688 4727 688
rect 4681 -700 4727 -688
rect 4777 688 4823 700
rect 4777 -688 4783 688
rect 4817 -688 4823 688
rect 4777 -700 4823 -688
rect 4873 688 4919 700
rect 4873 -688 4879 688
rect 4913 -688 4919 688
rect 4873 -700 4919 -688
rect 4969 688 5015 700
rect 4969 -688 4975 688
rect 5009 -688 5015 688
rect 4969 -700 5015 -688
rect 5065 688 5111 700
rect 5065 -688 5071 688
rect 5105 -688 5111 688
rect 5065 -700 5111 -688
rect 5161 688 5207 700
rect 5161 -688 5167 688
rect 5201 -688 5207 688
rect 5161 -700 5207 -688
rect 5257 688 5303 700
rect 5257 -688 5263 688
rect 5297 -688 5303 688
rect 5257 -700 5303 -688
rect 5353 688 5399 700
rect 5353 -688 5359 688
rect 5393 -688 5399 688
rect 5353 -700 5399 -688
rect 5449 688 5495 700
rect 5449 -688 5455 688
rect 5489 -688 5495 688
rect 5449 -700 5495 -688
rect 5545 688 5591 700
rect 5545 -688 5551 688
rect 5585 -688 5591 688
rect 5545 -700 5591 -688
rect 5641 688 5687 700
rect 5641 -688 5647 688
rect 5681 -688 5687 688
rect 5641 -700 5687 -688
rect 5737 688 5783 700
rect 5737 -688 5743 688
rect 5777 -688 5783 688
rect 5737 -700 5783 -688
rect 5833 688 5879 700
rect 5833 -688 5839 688
rect 5873 -688 5879 688
rect 5833 -700 5879 -688
rect 5929 688 5975 700
rect 5929 -688 5935 688
rect 5969 -688 5975 688
rect 5929 -700 5975 -688
rect 6025 688 6071 700
rect 6025 -688 6031 688
rect 6065 -688 6071 688
rect 6025 -700 6071 -688
rect 6121 688 6167 700
rect 6121 -688 6127 688
rect 6161 -688 6167 688
rect 6121 -700 6167 -688
rect 6217 688 6263 700
rect 6217 -688 6223 688
rect 6257 -688 6263 688
rect 6217 -700 6263 -688
rect 6313 688 6359 700
rect 6313 -688 6319 688
rect 6353 -688 6359 688
rect 6313 -700 6359 -688
rect 6409 688 6455 700
rect 6409 -688 6415 688
rect 6449 -688 6455 688
rect 6409 -700 6455 -688
rect 6505 688 6551 700
rect 6505 -688 6511 688
rect 6545 -688 6551 688
rect 6505 -700 6551 -688
rect 6601 688 6647 700
rect 6601 -688 6607 688
rect 6641 -688 6647 688
rect 6601 -700 6647 -688
rect 6697 688 6743 700
rect 6697 -688 6703 688
rect 6737 -688 6743 688
rect 6697 -700 6743 -688
rect 6793 688 6839 700
rect 6793 -688 6799 688
rect 6833 -688 6839 688
rect 6793 -700 6839 -688
rect 6889 688 6935 700
rect 6889 -688 6895 688
rect 6929 -688 6935 688
rect 6889 -700 6935 -688
rect 6985 688 7031 700
rect 6985 -688 6991 688
rect 7025 -688 7031 688
rect 6985 -700 7031 -688
rect 7081 688 7127 700
rect 7081 -688 7087 688
rect 7121 -688 7127 688
rect 7081 -700 7127 -688
rect 7177 688 7223 700
rect 7177 -688 7183 688
rect 7217 -688 7223 688
rect 7177 -700 7223 -688
rect 7273 688 7319 700
rect 7273 -688 7279 688
rect 7313 -688 7319 688
rect 7273 -700 7319 -688
rect 7369 688 7415 700
rect 7369 -688 7375 688
rect 7409 -688 7415 688
rect 7369 -700 7415 -688
rect 7465 688 7511 700
rect 7465 -688 7471 688
rect 7505 -688 7511 688
rect 7465 -700 7511 -688
rect 7561 688 7607 700
rect 7561 -688 7567 688
rect 7601 -688 7607 688
rect 7561 -700 7607 -688
rect 7657 688 7703 700
rect 7657 -688 7663 688
rect 7697 -688 7703 688
rect 7657 -700 7703 -688
rect 7753 688 7799 700
rect 7753 -688 7759 688
rect 7793 -688 7799 688
rect 7753 -700 7799 -688
rect 7849 688 7895 700
rect 7849 -688 7855 688
rect 7889 -688 7895 688
rect 7849 -700 7895 -688
rect 7945 688 7991 700
rect 7945 -688 7951 688
rect 7985 -688 7991 688
rect 7945 -700 7991 -688
rect 8041 688 8087 700
rect 8041 -688 8047 688
rect 8081 -688 8087 688
rect 8041 -700 8087 -688
rect 8137 688 8183 700
rect 8137 -688 8143 688
rect 8177 -688 8183 688
rect 8137 -700 8183 -688
rect 8233 688 8279 700
rect 8233 -688 8239 688
rect 8273 -688 8279 688
rect 8233 -700 8279 -688
rect 8329 688 8375 700
rect 8329 -688 8335 688
rect 8369 -688 8375 688
rect 8329 -700 8375 -688
rect 8425 688 8471 700
rect 8425 -688 8431 688
rect 8465 -688 8471 688
rect 8425 -700 8471 -688
rect 8521 688 8567 700
rect 8521 -688 8527 688
rect 8561 -688 8567 688
rect 8521 -700 8567 -688
rect 8617 688 8663 700
rect 8617 -688 8623 688
rect 8657 -688 8663 688
rect 8617 -700 8663 -688
rect 8713 688 8759 700
rect 8713 -688 8719 688
rect 8753 -688 8759 688
rect 8713 -700 8759 -688
rect 8809 688 8855 700
rect 8809 -688 8815 688
rect 8849 -688 8855 688
rect 8809 -700 8855 -688
rect 8905 688 8951 700
rect 8905 -688 8911 688
rect 8945 -688 8951 688
rect 8905 -700 8951 -688
rect 9001 688 9047 700
rect 9001 -688 9007 688
rect 9041 -688 9047 688
rect 9001 -700 9047 -688
rect 9097 688 9143 700
rect 9097 -688 9103 688
rect 9137 -688 9143 688
rect 9097 -700 9143 -688
rect 9193 688 9239 700
rect 9193 -688 9199 688
rect 9233 -688 9239 688
rect 9193 -700 9239 -688
rect 9289 688 9335 700
rect 9289 -688 9295 688
rect 9329 -688 9335 688
rect 9289 -700 9335 -688
rect 9385 688 9431 700
rect 9385 -688 9391 688
rect 9425 -688 9431 688
rect 9385 -700 9431 -688
rect 9481 688 9527 700
rect 9481 -688 9487 688
rect 9521 -688 9527 688
rect 9481 -700 9527 -688
rect 9577 688 9623 700
rect 9577 -688 9583 688
rect 9617 -688 9623 688
rect 9577 -700 9623 -688
rect 9673 688 9719 700
rect 9673 -688 9679 688
rect 9713 -688 9719 688
rect 9673 -700 9719 -688
rect 9769 688 9815 700
rect 9769 -688 9775 688
rect 9809 -688 9815 688
rect 9769 -700 9815 -688
rect 9865 688 9911 700
rect 9865 -688 9871 688
rect 9905 -688 9911 688
rect 9865 -700 9911 -688
rect 9961 688 10007 700
rect 9961 -688 9967 688
rect 10001 -688 10007 688
rect 9961 -700 10007 -688
rect 10057 688 10103 700
rect 10057 -688 10063 688
rect 10097 -688 10103 688
rect 10057 -700 10103 -688
rect 10153 688 10199 700
rect 10153 -688 10159 688
rect 10193 -688 10199 688
rect 10153 -700 10199 -688
rect 10249 688 10295 700
rect 10249 -688 10255 688
rect 10289 -688 10295 688
rect 10249 -700 10295 -688
rect 10345 688 10391 700
rect 10345 -688 10351 688
rect 10385 -688 10391 688
rect 10345 -700 10391 -688
rect 10441 688 10487 700
rect 10441 -688 10447 688
rect 10481 -688 10487 688
rect 10441 -700 10487 -688
rect 10537 688 10583 700
rect 10537 -688 10543 688
rect 10577 -688 10583 688
rect 10537 -700 10583 -688
rect -10541 -747 -10483 -741
rect -10541 -781 -10529 -747
rect -10495 -781 -10483 -747
rect -10541 -787 -10483 -781
rect -10349 -747 -10291 -741
rect -10349 -781 -10337 -747
rect -10303 -781 -10291 -747
rect -10349 -787 -10291 -781
rect -10157 -747 -10099 -741
rect -10157 -781 -10145 -747
rect -10111 -781 -10099 -747
rect -10157 -787 -10099 -781
rect -9965 -747 -9907 -741
rect -9965 -781 -9953 -747
rect -9919 -781 -9907 -747
rect -9965 -787 -9907 -781
rect -9773 -747 -9715 -741
rect -9773 -781 -9761 -747
rect -9727 -781 -9715 -747
rect -9773 -787 -9715 -781
rect -9581 -747 -9523 -741
rect -9581 -781 -9569 -747
rect -9535 -781 -9523 -747
rect -9581 -787 -9523 -781
rect -9389 -747 -9331 -741
rect -9389 -781 -9377 -747
rect -9343 -781 -9331 -747
rect -9389 -787 -9331 -781
rect -9197 -747 -9139 -741
rect -9197 -781 -9185 -747
rect -9151 -781 -9139 -747
rect -9197 -787 -9139 -781
rect -9005 -747 -8947 -741
rect -9005 -781 -8993 -747
rect -8959 -781 -8947 -747
rect -9005 -787 -8947 -781
rect -8813 -747 -8755 -741
rect -8813 -781 -8801 -747
rect -8767 -781 -8755 -747
rect -8813 -787 -8755 -781
rect -8621 -747 -8563 -741
rect -8621 -781 -8609 -747
rect -8575 -781 -8563 -747
rect -8621 -787 -8563 -781
rect -8429 -747 -8371 -741
rect -8429 -781 -8417 -747
rect -8383 -781 -8371 -747
rect -8429 -787 -8371 -781
rect -8237 -747 -8179 -741
rect -8237 -781 -8225 -747
rect -8191 -781 -8179 -747
rect -8237 -787 -8179 -781
rect -8045 -747 -7987 -741
rect -8045 -781 -8033 -747
rect -7999 -781 -7987 -747
rect -8045 -787 -7987 -781
rect -7853 -747 -7795 -741
rect -7853 -781 -7841 -747
rect -7807 -781 -7795 -747
rect -7853 -787 -7795 -781
rect -7661 -747 -7603 -741
rect -7661 -781 -7649 -747
rect -7615 -781 -7603 -747
rect -7661 -787 -7603 -781
rect -7469 -747 -7411 -741
rect -7469 -781 -7457 -747
rect -7423 -781 -7411 -747
rect -7469 -787 -7411 -781
rect -7277 -747 -7219 -741
rect -7277 -781 -7265 -747
rect -7231 -781 -7219 -747
rect -7277 -787 -7219 -781
rect -7085 -747 -7027 -741
rect -7085 -781 -7073 -747
rect -7039 -781 -7027 -747
rect -7085 -787 -7027 -781
rect -6893 -747 -6835 -741
rect -6893 -781 -6881 -747
rect -6847 -781 -6835 -747
rect -6893 -787 -6835 -781
rect -6701 -747 -6643 -741
rect -6701 -781 -6689 -747
rect -6655 -781 -6643 -747
rect -6701 -787 -6643 -781
rect -6509 -747 -6451 -741
rect -6509 -781 -6497 -747
rect -6463 -781 -6451 -747
rect -6509 -787 -6451 -781
rect -6317 -747 -6259 -741
rect -6317 -781 -6305 -747
rect -6271 -781 -6259 -747
rect -6317 -787 -6259 -781
rect -6125 -747 -6067 -741
rect -6125 -781 -6113 -747
rect -6079 -781 -6067 -747
rect -6125 -787 -6067 -781
rect -5933 -747 -5875 -741
rect -5933 -781 -5921 -747
rect -5887 -781 -5875 -747
rect -5933 -787 -5875 -781
rect -5741 -747 -5683 -741
rect -5741 -781 -5729 -747
rect -5695 -781 -5683 -747
rect -5741 -787 -5683 -781
rect -5549 -747 -5491 -741
rect -5549 -781 -5537 -747
rect -5503 -781 -5491 -747
rect -5549 -787 -5491 -781
rect -5357 -747 -5299 -741
rect -5357 -781 -5345 -747
rect -5311 -781 -5299 -747
rect -5357 -787 -5299 -781
rect -5165 -747 -5107 -741
rect -5165 -781 -5153 -747
rect -5119 -781 -5107 -747
rect -5165 -787 -5107 -781
rect -4973 -747 -4915 -741
rect -4973 -781 -4961 -747
rect -4927 -781 -4915 -747
rect -4973 -787 -4915 -781
rect -4781 -747 -4723 -741
rect -4781 -781 -4769 -747
rect -4735 -781 -4723 -747
rect -4781 -787 -4723 -781
rect -4589 -747 -4531 -741
rect -4589 -781 -4577 -747
rect -4543 -781 -4531 -747
rect -4589 -787 -4531 -781
rect -4397 -747 -4339 -741
rect -4397 -781 -4385 -747
rect -4351 -781 -4339 -747
rect -4397 -787 -4339 -781
rect -4205 -747 -4147 -741
rect -4205 -781 -4193 -747
rect -4159 -781 -4147 -747
rect -4205 -787 -4147 -781
rect -4013 -747 -3955 -741
rect -4013 -781 -4001 -747
rect -3967 -781 -3955 -747
rect -4013 -787 -3955 -781
rect -3821 -747 -3763 -741
rect -3821 -781 -3809 -747
rect -3775 -781 -3763 -747
rect -3821 -787 -3763 -781
rect -3629 -747 -3571 -741
rect -3629 -781 -3617 -747
rect -3583 -781 -3571 -747
rect -3629 -787 -3571 -781
rect -3437 -747 -3379 -741
rect -3437 -781 -3425 -747
rect -3391 -781 -3379 -747
rect -3437 -787 -3379 -781
rect -3245 -747 -3187 -741
rect -3245 -781 -3233 -747
rect -3199 -781 -3187 -747
rect -3245 -787 -3187 -781
rect -3053 -747 -2995 -741
rect -3053 -781 -3041 -747
rect -3007 -781 -2995 -747
rect -3053 -787 -2995 -781
rect -2861 -747 -2803 -741
rect -2861 -781 -2849 -747
rect -2815 -781 -2803 -747
rect -2861 -787 -2803 -781
rect -2669 -747 -2611 -741
rect -2669 -781 -2657 -747
rect -2623 -781 -2611 -747
rect -2669 -787 -2611 -781
rect -2477 -747 -2419 -741
rect -2477 -781 -2465 -747
rect -2431 -781 -2419 -747
rect -2477 -787 -2419 -781
rect -2285 -747 -2227 -741
rect -2285 -781 -2273 -747
rect -2239 -781 -2227 -747
rect -2285 -787 -2227 -781
rect -2093 -747 -2035 -741
rect -2093 -781 -2081 -747
rect -2047 -781 -2035 -747
rect -2093 -787 -2035 -781
rect -1901 -747 -1843 -741
rect -1901 -781 -1889 -747
rect -1855 -781 -1843 -747
rect -1901 -787 -1843 -781
rect -1709 -747 -1651 -741
rect -1709 -781 -1697 -747
rect -1663 -781 -1651 -747
rect -1709 -787 -1651 -781
rect -1517 -747 -1459 -741
rect -1517 -781 -1505 -747
rect -1471 -781 -1459 -747
rect -1517 -787 -1459 -781
rect -1325 -747 -1267 -741
rect -1325 -781 -1313 -747
rect -1279 -781 -1267 -747
rect -1325 -787 -1267 -781
rect -1133 -747 -1075 -741
rect -1133 -781 -1121 -747
rect -1087 -781 -1075 -747
rect -1133 -787 -1075 -781
rect -941 -747 -883 -741
rect -941 -781 -929 -747
rect -895 -781 -883 -747
rect -941 -787 -883 -781
rect -749 -747 -691 -741
rect -749 -781 -737 -747
rect -703 -781 -691 -747
rect -749 -787 -691 -781
rect -557 -747 -499 -741
rect -557 -781 -545 -747
rect -511 -781 -499 -747
rect -557 -787 -499 -781
rect -365 -747 -307 -741
rect -365 -781 -353 -747
rect -319 -781 -307 -747
rect -365 -787 -307 -781
rect -173 -747 -115 -741
rect -173 -781 -161 -747
rect -127 -781 -115 -747
rect -173 -787 -115 -781
rect 19 -747 77 -741
rect 19 -781 31 -747
rect 65 -781 77 -747
rect 19 -787 77 -781
rect 211 -747 269 -741
rect 211 -781 223 -747
rect 257 -781 269 -747
rect 211 -787 269 -781
rect 403 -747 461 -741
rect 403 -781 415 -747
rect 449 -781 461 -747
rect 403 -787 461 -781
rect 595 -747 653 -741
rect 595 -781 607 -747
rect 641 -781 653 -747
rect 595 -787 653 -781
rect 787 -747 845 -741
rect 787 -781 799 -747
rect 833 -781 845 -747
rect 787 -787 845 -781
rect 979 -747 1037 -741
rect 979 -781 991 -747
rect 1025 -781 1037 -747
rect 979 -787 1037 -781
rect 1171 -747 1229 -741
rect 1171 -781 1183 -747
rect 1217 -781 1229 -747
rect 1171 -787 1229 -781
rect 1363 -747 1421 -741
rect 1363 -781 1375 -747
rect 1409 -781 1421 -747
rect 1363 -787 1421 -781
rect 1555 -747 1613 -741
rect 1555 -781 1567 -747
rect 1601 -781 1613 -747
rect 1555 -787 1613 -781
rect 1747 -747 1805 -741
rect 1747 -781 1759 -747
rect 1793 -781 1805 -747
rect 1747 -787 1805 -781
rect 1939 -747 1997 -741
rect 1939 -781 1951 -747
rect 1985 -781 1997 -747
rect 1939 -787 1997 -781
rect 2131 -747 2189 -741
rect 2131 -781 2143 -747
rect 2177 -781 2189 -747
rect 2131 -787 2189 -781
rect 2323 -747 2381 -741
rect 2323 -781 2335 -747
rect 2369 -781 2381 -747
rect 2323 -787 2381 -781
rect 2515 -747 2573 -741
rect 2515 -781 2527 -747
rect 2561 -781 2573 -747
rect 2515 -787 2573 -781
rect 2707 -747 2765 -741
rect 2707 -781 2719 -747
rect 2753 -781 2765 -747
rect 2707 -787 2765 -781
rect 2899 -747 2957 -741
rect 2899 -781 2911 -747
rect 2945 -781 2957 -747
rect 2899 -787 2957 -781
rect 3091 -747 3149 -741
rect 3091 -781 3103 -747
rect 3137 -781 3149 -747
rect 3091 -787 3149 -781
rect 3283 -747 3341 -741
rect 3283 -781 3295 -747
rect 3329 -781 3341 -747
rect 3283 -787 3341 -781
rect 3475 -747 3533 -741
rect 3475 -781 3487 -747
rect 3521 -781 3533 -747
rect 3475 -787 3533 -781
rect 3667 -747 3725 -741
rect 3667 -781 3679 -747
rect 3713 -781 3725 -747
rect 3667 -787 3725 -781
rect 3859 -747 3917 -741
rect 3859 -781 3871 -747
rect 3905 -781 3917 -747
rect 3859 -787 3917 -781
rect 4051 -747 4109 -741
rect 4051 -781 4063 -747
rect 4097 -781 4109 -747
rect 4051 -787 4109 -781
rect 4243 -747 4301 -741
rect 4243 -781 4255 -747
rect 4289 -781 4301 -747
rect 4243 -787 4301 -781
rect 4435 -747 4493 -741
rect 4435 -781 4447 -747
rect 4481 -781 4493 -747
rect 4435 -787 4493 -781
rect 4627 -747 4685 -741
rect 4627 -781 4639 -747
rect 4673 -781 4685 -747
rect 4627 -787 4685 -781
rect 4819 -747 4877 -741
rect 4819 -781 4831 -747
rect 4865 -781 4877 -747
rect 4819 -787 4877 -781
rect 5011 -747 5069 -741
rect 5011 -781 5023 -747
rect 5057 -781 5069 -747
rect 5011 -787 5069 -781
rect 5203 -747 5261 -741
rect 5203 -781 5215 -747
rect 5249 -781 5261 -747
rect 5203 -787 5261 -781
rect 5395 -747 5453 -741
rect 5395 -781 5407 -747
rect 5441 -781 5453 -747
rect 5395 -787 5453 -781
rect 5587 -747 5645 -741
rect 5587 -781 5599 -747
rect 5633 -781 5645 -747
rect 5587 -787 5645 -781
rect 5779 -747 5837 -741
rect 5779 -781 5791 -747
rect 5825 -781 5837 -747
rect 5779 -787 5837 -781
rect 5971 -747 6029 -741
rect 5971 -781 5983 -747
rect 6017 -781 6029 -747
rect 5971 -787 6029 -781
rect 6163 -747 6221 -741
rect 6163 -781 6175 -747
rect 6209 -781 6221 -747
rect 6163 -787 6221 -781
rect 6355 -747 6413 -741
rect 6355 -781 6367 -747
rect 6401 -781 6413 -747
rect 6355 -787 6413 -781
rect 6547 -747 6605 -741
rect 6547 -781 6559 -747
rect 6593 -781 6605 -747
rect 6547 -787 6605 -781
rect 6739 -747 6797 -741
rect 6739 -781 6751 -747
rect 6785 -781 6797 -747
rect 6739 -787 6797 -781
rect 6931 -747 6989 -741
rect 6931 -781 6943 -747
rect 6977 -781 6989 -747
rect 6931 -787 6989 -781
rect 7123 -747 7181 -741
rect 7123 -781 7135 -747
rect 7169 -781 7181 -747
rect 7123 -787 7181 -781
rect 7315 -747 7373 -741
rect 7315 -781 7327 -747
rect 7361 -781 7373 -747
rect 7315 -787 7373 -781
rect 7507 -747 7565 -741
rect 7507 -781 7519 -747
rect 7553 -781 7565 -747
rect 7507 -787 7565 -781
rect 7699 -747 7757 -741
rect 7699 -781 7711 -747
rect 7745 -781 7757 -747
rect 7699 -787 7757 -781
rect 7891 -747 7949 -741
rect 7891 -781 7903 -747
rect 7937 -781 7949 -747
rect 7891 -787 7949 -781
rect 8083 -747 8141 -741
rect 8083 -781 8095 -747
rect 8129 -781 8141 -747
rect 8083 -787 8141 -781
rect 8275 -747 8333 -741
rect 8275 -781 8287 -747
rect 8321 -781 8333 -747
rect 8275 -787 8333 -781
rect 8467 -747 8525 -741
rect 8467 -781 8479 -747
rect 8513 -781 8525 -747
rect 8467 -787 8525 -781
rect 8659 -747 8717 -741
rect 8659 -781 8671 -747
rect 8705 -781 8717 -747
rect 8659 -787 8717 -781
rect 8851 -747 8909 -741
rect 8851 -781 8863 -747
rect 8897 -781 8909 -747
rect 8851 -787 8909 -781
rect 9043 -747 9101 -741
rect 9043 -781 9055 -747
rect 9089 -781 9101 -747
rect 9043 -787 9101 -781
rect 9235 -747 9293 -741
rect 9235 -781 9247 -747
rect 9281 -781 9293 -747
rect 9235 -787 9293 -781
rect 9427 -747 9485 -741
rect 9427 -781 9439 -747
rect 9473 -781 9485 -747
rect 9427 -787 9485 -781
rect 9619 -747 9677 -741
rect 9619 -781 9631 -747
rect 9665 -781 9677 -747
rect 9619 -787 9677 -781
rect 9811 -747 9869 -741
rect 9811 -781 9823 -747
rect 9857 -781 9869 -747
rect 9811 -787 9869 -781
rect 10003 -747 10061 -741
rect 10003 -781 10015 -747
rect 10049 -781 10061 -747
rect 10003 -787 10061 -781
rect 10195 -747 10253 -741
rect 10195 -781 10207 -747
rect 10241 -781 10253 -747
rect 10195 -787 10253 -781
rect 10387 -747 10445 -741
rect 10387 -781 10399 -747
rect 10433 -781 10445 -747
rect 10387 -787 10445 -781
<< properties >>
string FIXED_BBOX -10674 -866 10674 866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 0.15 m 1 nf 220 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
