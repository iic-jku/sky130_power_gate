magic
tech sky130A
magscale 1 2
timestamp 1697723814
<< viali >>
rect 328 21868 882 21932
<< metal1 >>
rect 122 22286 1716 22304
rect 122 22222 132 22286
rect 1706 22222 1716 22286
rect 122 22204 1716 22222
rect 132 828 178 22204
rect 316 21934 894 21938
rect 316 21932 352 21934
rect 858 21932 894 21934
rect 316 21868 328 21932
rect 882 21868 894 21932
rect 316 21862 894 21868
rect 1660 732 1706 22204
<< via1 >>
rect 132 22222 1706 22286
rect 352 21932 858 21934
rect 342 21868 868 21932
<< metal2 >>
rect 132 22286 1706 22296
rect 132 22212 1706 22222
rect 342 21934 868 21942
rect 342 21932 352 21934
rect 858 21932 868 21934
rect 342 21858 868 21868
<< via2 >>
rect 132 22222 1706 22286
rect 352 21868 858 21934
<< metal3 >>
rect 122 22286 1716 22291
rect 122 22222 132 22286
rect 1706 22222 1716 22286
rect 122 22217 1716 22222
rect 344 21934 868 21944
rect 344 21868 352 21934
rect 858 21868 868 21934
rect 344 21820 868 21868
<< via3 >>
rect 132 22222 1706 22286
rect 352 21868 858 21934
<< metal4 >>
rect 0 22286 1840 22304
rect 0 22222 132 22286
rect 1706 22222 1840 22286
rect 0 22204 1840 22222
rect 0 0 240 22000
rect 340 21934 870 22000
rect 340 21868 352 21934
rect 858 21868 870 21934
rect 340 2089 870 21868
rect 339 2023 871 2089
rect 340 1899 870 2023
rect 339 1833 871 1899
rect 340 1705 870 1833
rect 339 1639 871 1705
rect 340 1515 870 1639
rect 339 1449 871 1515
rect 340 1323 870 1449
rect 339 1257 871 1323
rect 340 1129 870 1257
rect 339 1063 871 1129
rect 340 939 870 1063
rect 339 873 871 939
rect 340 747 870 873
rect 339 681 871 747
rect 340 0 870 681
rect 970 0 1500 22000
rect 1600 0 1840 22000
use cont_even  cont_even_0
timestamp 1697722671
transform 0 1 918 -1 0 11217
box -10603 -576 10603 -50
use cont_odd  cont_odd_0
timestamp 1697723018
transform 0 1 918 -1 0 11217
box -10507 52 10507 582
use sky130_fd_pr__pfet_01v8_6QHARF  sky130_fd_pr__pfet_01v8_6QHARF_0
timestamp 1697193002
transform 0 1 919 -1 0 11217
box -10727 -919 10727 919
<< labels >>
rlabel metal4 0 0 240 22000 1 VGND
port 1 n ground input
rlabel metal4 1600 0 1840 22000 1 VGND
port 1 n ground input
rlabel metal4 340 0 870 22000 1 VPWR
port 2 n power input
rlabel metal4 970 0 1500 22000 1 GPWR
port 3 n power output
rlabel metal4 0 22204 1840 22304 1 ctrl
port 4 n signal input
<< end >>
