magic
tech sky130A
magscale 1 2
timestamp 1697796922
<< error_s >>
rect 339 2044 399 2089
rect 339 2023 400 2044
rect 342 1963 400 2023
rect 810 1963 868 2044
rect 870 2023 930 2089
rect 342 1958 400 1959
rect 810 1958 868 1959
rect 339 1852 399 1899
rect 339 1833 400 1852
rect 342 1773 400 1833
rect 810 1773 868 1852
rect 870 1833 930 1899
rect 339 1660 399 1705
rect 339 1639 400 1660
rect 342 1579 400 1639
rect 810 1579 868 1660
rect 870 1639 930 1705
rect 342 1574 400 1575
rect 810 1574 868 1575
rect 339 1468 399 1515
rect 339 1449 400 1468
rect 342 1389 400 1449
rect 810 1389 868 1468
rect 870 1449 930 1515
rect 342 1382 400 1383
rect 810 1382 868 1383
rect 339 1276 399 1323
rect 339 1257 400 1276
rect 342 1197 400 1257
rect 810 1197 868 1276
rect 870 1257 930 1323
rect 339 1084 399 1129
rect 339 1063 400 1084
rect 342 1003 400 1063
rect 810 1003 868 1084
rect 870 1063 930 1129
rect 342 998 400 999
rect 810 998 868 999
rect 339 892 399 939
rect 339 873 400 892
rect 342 813 400 873
rect 810 813 868 892
rect 870 873 930 939
rect 342 806 400 807
rect 810 806 868 807
rect 339 700 399 747
rect 339 681 400 700
rect 342 621 400 681
rect 810 621 868 700
rect 870 681 930 747
<< metal1 >>
rect 132 828 178 21710
rect 1660 732 1706 21844
<< metal4 >>
rect 339 2023 340 2089
rect 870 2023 871 2089
rect 339 1833 340 1899
rect 870 1833 871 1899
rect 339 1639 340 1705
rect 870 1639 871 1705
rect 339 1449 340 1515
rect 870 1449 871 1515
rect 339 1257 340 1323
rect 870 1257 871 1323
rect 339 1063 340 1129
rect 870 1063 871 1129
rect 339 873 340 939
rect 870 873 871 939
rect 339 681 340 747
rect 870 681 871 747
use cont_even  cont_even_0
timestamp 1697722671
transform 0 1 918 -1 0 11217
box -10603 -576 10603 -50
use cont_odd  cont_odd_0
timestamp 1697723018
transform 0 1 918 -1 0 11217
box -10507 52 10507 582
use sky130_fd_pr__pfet_01v8_6QHARF  sky130_fd_pr__pfet_01v8_6QHARF_0
timestamp 1697193002
transform 0 1 919 -1 0 11217
box -10727 -919 10727 919
<< end >>
