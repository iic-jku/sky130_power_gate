magic
tech sky130A
magscale 1 2
timestamp 1697723018
<< metal1 >>
rect -10497 572 -10431 582
rect -10497 52 -10431 62
rect -10305 572 -10239 582
rect -10305 52 -10239 62
rect -10113 572 -10047 582
rect -10113 52 -10047 62
rect -9921 572 -9855 582
rect -9921 52 -9855 62
rect -9729 572 -9663 582
rect -9729 52 -9663 62
rect -9537 572 -9471 582
rect -9537 52 -9471 62
rect -9345 572 -9279 582
rect -9345 52 -9279 62
rect -9153 572 -9087 582
rect -9153 52 -9087 62
rect -8961 572 -8895 582
rect -8961 52 -8895 62
rect -8769 572 -8703 582
rect -8769 52 -8703 62
rect -8577 572 -8511 582
rect -8577 52 -8511 62
rect -8385 572 -8319 582
rect -8385 52 -8319 62
rect -8193 572 -8127 582
rect -8193 52 -8127 62
rect -8001 572 -7935 582
rect -8001 52 -7935 62
rect -7809 572 -7743 582
rect -7809 52 -7743 62
rect -7617 572 -7551 582
rect -7617 52 -7551 62
rect -7425 572 -7359 582
rect -7425 52 -7359 62
rect -7233 572 -7167 582
rect -7233 52 -7167 62
rect -7041 572 -6975 582
rect -7041 52 -6975 62
rect -6849 572 -6783 582
rect -6849 52 -6783 62
rect -6657 572 -6591 582
rect -6657 52 -6591 62
rect -6465 572 -6399 582
rect -6465 52 -6399 62
rect -6273 572 -6207 582
rect -6273 52 -6207 62
rect -6081 572 -6015 582
rect -6081 52 -6015 62
rect -5889 572 -5823 582
rect -5889 52 -5823 62
rect -5697 572 -5631 582
rect -5697 52 -5631 62
rect -5505 572 -5439 582
rect -5505 52 -5439 62
rect -5313 572 -5247 582
rect -5313 52 -5247 62
rect -5121 572 -5055 582
rect -5121 52 -5055 62
rect -4929 572 -4863 582
rect -4929 52 -4863 62
rect -4737 572 -4671 582
rect -4737 52 -4671 62
rect -4545 572 -4479 582
rect -4545 52 -4479 62
rect -4353 572 -4287 582
rect -4353 52 -4287 62
rect -4161 572 -4095 582
rect -4161 52 -4095 62
rect -3969 572 -3903 582
rect -3969 52 -3903 62
rect -3777 572 -3711 582
rect -3777 52 -3711 62
rect -3585 572 -3519 582
rect -3585 52 -3519 62
rect -3393 572 -3327 582
rect -3393 52 -3327 62
rect -3201 572 -3135 582
rect -3201 52 -3135 62
rect -3009 572 -2943 582
rect -3009 52 -2943 62
rect -2817 572 -2751 582
rect -2817 52 -2751 62
rect -2625 572 -2559 582
rect -2625 52 -2559 62
rect -2433 572 -2367 582
rect -2433 52 -2367 62
rect -2241 572 -2175 582
rect -2241 52 -2175 62
rect -2049 572 -1983 582
rect -2049 52 -1983 62
rect -1857 572 -1791 582
rect -1857 52 -1791 62
rect -1665 572 -1599 582
rect -1665 52 -1599 62
rect -1473 572 -1407 582
rect -1473 52 -1407 62
rect -1281 572 -1215 582
rect -1281 52 -1215 62
rect -1089 572 -1023 582
rect -1089 52 -1023 62
rect -897 572 -831 582
rect -897 52 -831 62
rect -705 572 -639 582
rect -705 52 -639 62
rect -513 572 -447 582
rect -513 52 -447 62
rect -321 572 -255 582
rect -321 52 -255 62
rect -129 572 -63 582
rect -129 52 -63 62
rect 63 572 129 582
rect 63 52 129 62
rect 255 572 321 582
rect 255 52 321 62
rect 447 572 513 582
rect 447 52 513 62
rect 639 572 705 582
rect 639 52 705 62
rect 831 572 897 582
rect 831 52 897 62
rect 1023 572 1089 582
rect 1023 52 1089 62
rect 1215 572 1281 582
rect 1215 52 1281 62
rect 1407 572 1473 582
rect 1407 52 1473 62
rect 1599 572 1665 582
rect 1599 52 1665 62
rect 1791 572 1857 582
rect 1791 52 1857 62
rect 1983 572 2049 582
rect 1983 52 2049 62
rect 2175 572 2241 582
rect 2175 52 2241 62
rect 2367 572 2433 582
rect 2367 52 2433 62
rect 2559 572 2625 582
rect 2559 52 2625 62
rect 2751 572 2817 582
rect 2751 52 2817 62
rect 2943 572 3009 582
rect 2943 52 3009 62
rect 3135 572 3201 582
rect 3135 52 3201 62
rect 3327 572 3393 582
rect 3327 52 3393 62
rect 3519 572 3585 582
rect 3519 52 3585 62
rect 3711 572 3777 582
rect 3711 52 3777 62
rect 3903 572 3969 582
rect 3903 52 3969 62
rect 4095 572 4161 582
rect 4095 52 4161 62
rect 4287 572 4353 582
rect 4287 52 4353 62
rect 4479 572 4545 582
rect 4479 52 4545 62
rect 4671 572 4737 582
rect 4671 52 4737 62
rect 4863 572 4929 582
rect 4863 52 4929 62
rect 5055 572 5121 582
rect 5055 52 5121 62
rect 5247 572 5313 582
rect 5247 52 5313 62
rect 5439 572 5505 582
rect 5439 52 5505 62
rect 5631 572 5697 582
rect 5631 52 5697 62
rect 5823 572 5889 582
rect 5823 52 5889 62
rect 6015 572 6081 582
rect 6015 52 6081 62
rect 6207 572 6273 582
rect 6207 52 6273 62
rect 6399 572 6465 582
rect 6399 52 6465 62
rect 6591 572 6657 582
rect 6591 52 6657 62
rect 6783 572 6849 582
rect 6783 52 6849 62
rect 6975 572 7041 582
rect 6975 52 7041 62
rect 7167 572 7233 582
rect 7167 52 7233 62
rect 7359 572 7425 582
rect 7359 52 7425 62
rect 7551 572 7617 582
rect 7551 52 7617 62
rect 7743 572 7809 582
rect 7743 52 7809 62
rect 7935 572 8001 582
rect 7935 52 8001 62
rect 8127 572 8193 582
rect 8127 52 8193 62
rect 8319 572 8385 582
rect 8319 52 8385 62
rect 8511 572 8577 582
rect 8511 52 8577 62
rect 8703 572 8769 582
rect 8703 52 8769 62
rect 8895 572 8961 582
rect 8895 52 8961 62
rect 9087 572 9153 582
rect 9087 52 9153 62
rect 9279 572 9345 582
rect 9279 52 9345 62
rect 9471 572 9537 582
rect 9471 52 9537 62
rect 9663 572 9729 582
rect 9663 52 9729 62
rect 9855 572 9921 582
rect 9855 52 9921 62
rect 10047 572 10113 582
rect 10047 52 10113 62
rect 10239 572 10305 582
rect 10239 52 10305 62
rect 10431 572 10497 582
rect 10431 52 10497 62
<< via1 >>
rect -10497 62 -10431 572
rect -10305 62 -10239 572
rect -10113 62 -10047 572
rect -9921 62 -9855 572
rect -9729 62 -9663 572
rect -9537 62 -9471 572
rect -9345 62 -9279 572
rect -9153 62 -9087 572
rect -8961 62 -8895 572
rect -8769 62 -8703 572
rect -8577 62 -8511 572
rect -8385 62 -8319 572
rect -8193 62 -8127 572
rect -8001 62 -7935 572
rect -7809 62 -7743 572
rect -7617 62 -7551 572
rect -7425 62 -7359 572
rect -7233 62 -7167 572
rect -7041 62 -6975 572
rect -6849 62 -6783 572
rect -6657 62 -6591 572
rect -6465 62 -6399 572
rect -6273 62 -6207 572
rect -6081 62 -6015 572
rect -5889 62 -5823 572
rect -5697 62 -5631 572
rect -5505 62 -5439 572
rect -5313 62 -5247 572
rect -5121 62 -5055 572
rect -4929 62 -4863 572
rect -4737 62 -4671 572
rect -4545 62 -4479 572
rect -4353 62 -4287 572
rect -4161 62 -4095 572
rect -3969 62 -3903 572
rect -3777 62 -3711 572
rect -3585 62 -3519 572
rect -3393 62 -3327 572
rect -3201 62 -3135 572
rect -3009 62 -2943 572
rect -2817 62 -2751 572
rect -2625 62 -2559 572
rect -2433 62 -2367 572
rect -2241 62 -2175 572
rect -2049 62 -1983 572
rect -1857 62 -1791 572
rect -1665 62 -1599 572
rect -1473 62 -1407 572
rect -1281 62 -1215 572
rect -1089 62 -1023 572
rect -897 62 -831 572
rect -705 62 -639 572
rect -513 62 -447 572
rect -321 62 -255 572
rect -129 62 -63 572
rect 63 62 129 572
rect 255 62 321 572
rect 447 62 513 572
rect 639 62 705 572
rect 831 62 897 572
rect 1023 62 1089 572
rect 1215 62 1281 572
rect 1407 62 1473 572
rect 1599 62 1665 572
rect 1791 62 1857 572
rect 1983 62 2049 572
rect 2175 62 2241 572
rect 2367 62 2433 572
rect 2559 62 2625 572
rect 2751 62 2817 572
rect 2943 62 3009 572
rect 3135 62 3201 572
rect 3327 62 3393 572
rect 3519 62 3585 572
rect 3711 62 3777 572
rect 3903 62 3969 572
rect 4095 62 4161 572
rect 4287 62 4353 572
rect 4479 62 4545 572
rect 4671 62 4737 572
rect 4863 62 4929 572
rect 5055 62 5121 572
rect 5247 62 5313 572
rect 5439 62 5505 572
rect 5631 62 5697 572
rect 5823 62 5889 572
rect 6015 62 6081 572
rect 6207 62 6273 572
rect 6399 62 6465 572
rect 6591 62 6657 572
rect 6783 62 6849 572
rect 6975 62 7041 572
rect 7167 62 7233 572
rect 7359 62 7425 572
rect 7551 62 7617 572
rect 7743 62 7809 572
rect 7935 62 8001 572
rect 8127 62 8193 572
rect 8319 62 8385 572
rect 8511 62 8577 572
rect 8703 62 8769 572
rect 8895 62 8961 572
rect 9087 62 9153 572
rect 9279 62 9345 572
rect 9471 62 9537 572
rect 9663 62 9729 572
rect 9855 62 9921 572
rect 10047 62 10113 572
rect 10239 62 10305 572
rect 10431 62 10497 572
<< metal2 >>
rect -10507 572 -10421 582
rect -10507 62 -10497 572
rect -10431 62 -10421 572
rect -10507 52 -10421 62
rect -10315 572 -10229 582
rect -10315 62 -10305 572
rect -10239 62 -10229 572
rect -10315 52 -10229 62
rect -10123 572 -10037 582
rect -10123 62 -10113 572
rect -10047 62 -10037 572
rect -10123 52 -10037 62
rect -9931 572 -9845 582
rect -9931 62 -9921 572
rect -9855 62 -9845 572
rect -9931 52 -9845 62
rect -9739 572 -9653 582
rect -9739 62 -9729 572
rect -9663 62 -9653 572
rect -9739 52 -9653 62
rect -9547 572 -9461 582
rect -9547 62 -9537 572
rect -9471 62 -9461 572
rect -9547 52 -9461 62
rect -9355 572 -9269 582
rect -9355 62 -9345 572
rect -9279 62 -9269 572
rect -9355 52 -9269 62
rect -9163 572 -9077 582
rect -9163 62 -9153 572
rect -9087 62 -9077 572
rect -9163 52 -9077 62
rect -8971 572 -8885 582
rect -8971 62 -8961 572
rect -8895 62 -8885 572
rect -8971 52 -8885 62
rect -8779 572 -8693 582
rect -8779 62 -8769 572
rect -8703 62 -8693 572
rect -8779 52 -8693 62
rect -8587 572 -8501 582
rect -8587 62 -8577 572
rect -8511 62 -8501 572
rect -8587 52 -8501 62
rect -8395 572 -8309 582
rect -8395 62 -8385 572
rect -8319 62 -8309 572
rect -8395 52 -8309 62
rect -8203 572 -8117 582
rect -8203 62 -8193 572
rect -8127 62 -8117 572
rect -8203 52 -8117 62
rect -8011 572 -7925 582
rect -8011 62 -8001 572
rect -7935 62 -7925 572
rect -8011 52 -7925 62
rect -7819 572 -7733 582
rect -7819 62 -7809 572
rect -7743 62 -7733 572
rect -7819 52 -7733 62
rect -7627 572 -7541 582
rect -7627 62 -7617 572
rect -7551 62 -7541 572
rect -7627 52 -7541 62
rect -7435 572 -7349 582
rect -7435 62 -7425 572
rect -7359 62 -7349 572
rect -7435 52 -7349 62
rect -7243 572 -7157 582
rect -7243 62 -7233 572
rect -7167 62 -7157 572
rect -7243 52 -7157 62
rect -7051 572 -6965 582
rect -7051 62 -7041 572
rect -6975 62 -6965 572
rect -7051 52 -6965 62
rect -6859 572 -6773 582
rect -6859 62 -6849 572
rect -6783 62 -6773 572
rect -6859 52 -6773 62
rect -6667 572 -6581 582
rect -6667 62 -6657 572
rect -6591 62 -6581 572
rect -6667 52 -6581 62
rect -6475 572 -6389 582
rect -6475 62 -6465 572
rect -6399 62 -6389 572
rect -6475 52 -6389 62
rect -6283 572 -6197 582
rect -6283 62 -6273 572
rect -6207 62 -6197 572
rect -6283 52 -6197 62
rect -6091 572 -6005 582
rect -6091 62 -6081 572
rect -6015 62 -6005 572
rect -6091 52 -6005 62
rect -5899 572 -5813 582
rect -5899 62 -5889 572
rect -5823 62 -5813 572
rect -5899 52 -5813 62
rect -5707 572 -5621 582
rect -5707 62 -5697 572
rect -5631 62 -5621 572
rect -5707 52 -5621 62
rect -5515 572 -5429 582
rect -5515 62 -5505 572
rect -5439 62 -5429 572
rect -5515 52 -5429 62
rect -5323 572 -5237 582
rect -5323 62 -5313 572
rect -5247 62 -5237 572
rect -5323 52 -5237 62
rect -5131 572 -5045 582
rect -5131 62 -5121 572
rect -5055 62 -5045 572
rect -5131 52 -5045 62
rect -4939 572 -4853 582
rect -4939 62 -4929 572
rect -4863 62 -4853 572
rect -4939 52 -4853 62
rect -4747 572 -4661 582
rect -4747 62 -4737 572
rect -4671 62 -4661 572
rect -4747 52 -4661 62
rect -4555 572 -4469 582
rect -4555 62 -4545 572
rect -4479 62 -4469 572
rect -4555 52 -4469 62
rect -4363 572 -4277 582
rect -4363 62 -4353 572
rect -4287 62 -4277 572
rect -4363 52 -4277 62
rect -4171 572 -4085 582
rect -4171 62 -4161 572
rect -4095 62 -4085 572
rect -4171 52 -4085 62
rect -3979 572 -3893 582
rect -3979 62 -3969 572
rect -3903 62 -3893 572
rect -3979 52 -3893 62
rect -3787 572 -3701 582
rect -3787 62 -3777 572
rect -3711 62 -3701 572
rect -3787 52 -3701 62
rect -3595 572 -3509 582
rect -3595 62 -3585 572
rect -3519 62 -3509 572
rect -3595 52 -3509 62
rect -3403 572 -3317 582
rect -3403 62 -3393 572
rect -3327 62 -3317 572
rect -3403 52 -3317 62
rect -3211 572 -3125 582
rect -3211 62 -3201 572
rect -3135 62 -3125 572
rect -3211 52 -3125 62
rect -3019 572 -2933 582
rect -3019 62 -3009 572
rect -2943 62 -2933 572
rect -3019 52 -2933 62
rect -2827 572 -2741 582
rect -2827 62 -2817 572
rect -2751 62 -2741 572
rect -2827 52 -2741 62
rect -2635 572 -2549 582
rect -2635 62 -2625 572
rect -2559 62 -2549 572
rect -2635 52 -2549 62
rect -2443 572 -2357 582
rect -2443 62 -2433 572
rect -2367 62 -2357 572
rect -2443 52 -2357 62
rect -2251 572 -2165 582
rect -2251 62 -2241 572
rect -2175 62 -2165 572
rect -2251 52 -2165 62
rect -2059 572 -1973 582
rect -2059 62 -2049 572
rect -1983 62 -1973 572
rect -2059 52 -1973 62
rect -1867 572 -1781 582
rect -1867 62 -1857 572
rect -1791 62 -1781 572
rect -1867 52 -1781 62
rect -1675 572 -1589 582
rect -1675 62 -1665 572
rect -1599 62 -1589 572
rect -1675 52 -1589 62
rect -1483 572 -1397 582
rect -1483 62 -1473 572
rect -1407 62 -1397 572
rect -1483 52 -1397 62
rect -1291 572 -1205 582
rect -1291 62 -1281 572
rect -1215 62 -1205 572
rect -1291 52 -1205 62
rect -1099 572 -1013 582
rect -1099 62 -1089 572
rect -1023 62 -1013 572
rect -1099 52 -1013 62
rect -907 572 -821 582
rect -907 62 -897 572
rect -831 62 -821 572
rect -907 52 -821 62
rect -715 572 -629 582
rect -715 62 -705 572
rect -639 62 -629 572
rect -715 52 -629 62
rect -523 572 -437 582
rect -523 62 -513 572
rect -447 62 -437 572
rect -523 52 -437 62
rect -331 572 -245 582
rect -331 62 -321 572
rect -255 62 -245 572
rect -331 52 -245 62
rect -139 572 -53 582
rect -139 62 -129 572
rect -63 62 -53 572
rect -139 52 -53 62
rect 53 572 139 582
rect 53 62 63 572
rect 129 62 139 572
rect 53 52 139 62
rect 245 572 331 582
rect 245 62 255 572
rect 321 62 331 572
rect 245 52 331 62
rect 437 572 523 582
rect 437 62 447 572
rect 513 62 523 572
rect 437 52 523 62
rect 629 572 715 582
rect 629 62 639 572
rect 705 62 715 572
rect 629 52 715 62
rect 821 572 907 582
rect 821 62 831 572
rect 897 62 907 572
rect 821 52 907 62
rect 1013 572 1099 582
rect 1013 62 1023 572
rect 1089 62 1099 572
rect 1013 52 1099 62
rect 1205 572 1291 582
rect 1205 62 1215 572
rect 1281 62 1291 572
rect 1205 52 1291 62
rect 1397 572 1483 582
rect 1397 62 1407 572
rect 1473 62 1483 572
rect 1397 52 1483 62
rect 1589 572 1675 582
rect 1589 62 1599 572
rect 1665 62 1675 572
rect 1589 52 1675 62
rect 1781 572 1867 582
rect 1781 62 1791 572
rect 1857 62 1867 572
rect 1781 52 1867 62
rect 1973 572 2059 582
rect 1973 62 1983 572
rect 2049 62 2059 572
rect 1973 52 2059 62
rect 2165 572 2251 582
rect 2165 62 2175 572
rect 2241 62 2251 572
rect 2165 52 2251 62
rect 2357 572 2443 582
rect 2357 62 2367 572
rect 2433 62 2443 572
rect 2357 52 2443 62
rect 2549 572 2635 582
rect 2549 62 2559 572
rect 2625 62 2635 572
rect 2549 52 2635 62
rect 2741 572 2827 582
rect 2741 62 2751 572
rect 2817 62 2827 572
rect 2741 52 2827 62
rect 2933 572 3019 582
rect 2933 62 2943 572
rect 3009 62 3019 572
rect 2933 52 3019 62
rect 3125 572 3211 582
rect 3125 62 3135 572
rect 3201 62 3211 572
rect 3125 52 3211 62
rect 3317 572 3403 582
rect 3317 62 3327 572
rect 3393 62 3403 572
rect 3317 52 3403 62
rect 3509 572 3595 582
rect 3509 62 3519 572
rect 3585 62 3595 572
rect 3509 52 3595 62
rect 3701 572 3787 582
rect 3701 62 3711 572
rect 3777 62 3787 572
rect 3701 52 3787 62
rect 3893 572 3979 582
rect 3893 62 3903 572
rect 3969 62 3979 572
rect 3893 52 3979 62
rect 4085 572 4171 582
rect 4085 62 4095 572
rect 4161 62 4171 572
rect 4085 52 4171 62
rect 4277 572 4363 582
rect 4277 62 4287 572
rect 4353 62 4363 572
rect 4277 52 4363 62
rect 4469 572 4555 582
rect 4469 62 4479 572
rect 4545 62 4555 572
rect 4469 52 4555 62
rect 4661 572 4747 582
rect 4661 62 4671 572
rect 4737 62 4747 572
rect 4661 52 4747 62
rect 4853 572 4939 582
rect 4853 62 4863 572
rect 4929 62 4939 572
rect 4853 52 4939 62
rect 5045 572 5131 582
rect 5045 62 5055 572
rect 5121 62 5131 572
rect 5045 52 5131 62
rect 5237 572 5323 582
rect 5237 62 5247 572
rect 5313 62 5323 572
rect 5237 52 5323 62
rect 5429 572 5515 582
rect 5429 62 5439 572
rect 5505 62 5515 572
rect 5429 52 5515 62
rect 5621 572 5707 582
rect 5621 62 5631 572
rect 5697 62 5707 572
rect 5621 52 5707 62
rect 5813 572 5899 582
rect 5813 62 5823 572
rect 5889 62 5899 572
rect 5813 52 5899 62
rect 6005 572 6091 582
rect 6005 62 6015 572
rect 6081 62 6091 572
rect 6005 52 6091 62
rect 6197 572 6283 582
rect 6197 62 6207 572
rect 6273 62 6283 572
rect 6197 52 6283 62
rect 6389 572 6475 582
rect 6389 62 6399 572
rect 6465 62 6475 572
rect 6389 52 6475 62
rect 6581 572 6667 582
rect 6581 62 6591 572
rect 6657 62 6667 572
rect 6581 52 6667 62
rect 6773 572 6859 582
rect 6773 62 6783 572
rect 6849 62 6859 572
rect 6773 52 6859 62
rect 6965 572 7051 582
rect 6965 62 6975 572
rect 7041 62 7051 572
rect 6965 52 7051 62
rect 7157 572 7243 582
rect 7157 62 7167 572
rect 7233 62 7243 572
rect 7157 52 7243 62
rect 7349 572 7435 582
rect 7349 62 7359 572
rect 7425 62 7435 572
rect 7349 52 7435 62
rect 7541 572 7627 582
rect 7541 62 7551 572
rect 7617 62 7627 572
rect 7541 52 7627 62
rect 7733 572 7819 582
rect 7733 62 7743 572
rect 7809 62 7819 572
rect 7733 52 7819 62
rect 7925 572 8011 582
rect 7925 62 7935 572
rect 8001 62 8011 572
rect 7925 52 8011 62
rect 8117 572 8203 582
rect 8117 62 8127 572
rect 8193 62 8203 572
rect 8117 52 8203 62
rect 8309 572 8395 582
rect 8309 62 8319 572
rect 8385 62 8395 572
rect 8309 52 8395 62
rect 8501 572 8587 582
rect 8501 62 8511 572
rect 8577 62 8587 572
rect 8501 52 8587 62
rect 8693 572 8779 582
rect 8693 62 8703 572
rect 8769 62 8779 572
rect 8693 52 8779 62
rect 8885 572 8971 582
rect 8885 62 8895 572
rect 8961 62 8971 572
rect 8885 52 8971 62
rect 9077 572 9163 582
rect 9077 62 9087 572
rect 9153 62 9163 572
rect 9077 52 9163 62
rect 9269 572 9355 582
rect 9269 62 9279 572
rect 9345 62 9355 572
rect 9269 52 9355 62
rect 9461 572 9547 582
rect 9461 62 9471 572
rect 9537 62 9547 572
rect 9461 52 9547 62
rect 9653 572 9739 582
rect 9653 62 9663 572
rect 9729 62 9739 572
rect 9653 52 9739 62
rect 9845 572 9931 582
rect 9845 62 9855 572
rect 9921 62 9931 572
rect 9845 52 9931 62
rect 10037 572 10123 582
rect 10037 62 10047 572
rect 10113 62 10123 572
rect 10037 52 10123 62
rect 10229 572 10315 582
rect 10229 62 10239 572
rect 10305 62 10315 572
rect 10229 52 10315 62
rect 10421 572 10507 582
rect 10421 62 10431 572
rect 10497 62 10507 572
rect 10421 52 10507 62
<< via2 >>
rect -10497 62 -10431 572
rect -10305 62 -10239 572
rect -10113 62 -10047 572
rect -9921 62 -9855 572
rect -9729 62 -9663 572
rect -9537 62 -9471 572
rect -9345 62 -9279 572
rect -9153 62 -9087 572
rect -8961 62 -8895 572
rect -8769 62 -8703 572
rect -8577 62 -8511 572
rect -8385 62 -8319 572
rect -8193 62 -8127 572
rect -8001 62 -7935 572
rect -7809 62 -7743 572
rect -7617 62 -7551 572
rect -7425 62 -7359 572
rect -7233 62 -7167 572
rect -7041 62 -6975 572
rect -6849 62 -6783 572
rect -6657 62 -6591 572
rect -6465 62 -6399 572
rect -6273 62 -6207 572
rect -6081 62 -6015 572
rect -5889 62 -5823 572
rect -5697 62 -5631 572
rect -5505 62 -5439 572
rect -5313 62 -5247 572
rect -5121 62 -5055 572
rect -4929 62 -4863 572
rect -4737 62 -4671 572
rect -4545 62 -4479 572
rect -4353 62 -4287 572
rect -4161 62 -4095 572
rect -3969 62 -3903 572
rect -3777 62 -3711 572
rect -3585 62 -3519 572
rect -3393 62 -3327 572
rect -3201 62 -3135 572
rect -3009 62 -2943 572
rect -2817 62 -2751 572
rect -2625 62 -2559 572
rect -2433 62 -2367 572
rect -2241 62 -2175 572
rect -2049 62 -1983 572
rect -1857 62 -1791 572
rect -1665 62 -1599 572
rect -1473 62 -1407 572
rect -1281 62 -1215 572
rect -1089 62 -1023 572
rect -897 62 -831 572
rect -705 62 -639 572
rect -513 62 -447 572
rect -321 62 -255 572
rect -129 62 -63 572
rect 63 62 129 572
rect 255 62 321 572
rect 447 62 513 572
rect 639 62 705 572
rect 831 62 897 572
rect 1023 62 1089 572
rect 1215 62 1281 572
rect 1407 62 1473 572
rect 1599 62 1665 572
rect 1791 62 1857 572
rect 1983 62 2049 572
rect 2175 62 2241 572
rect 2367 62 2433 572
rect 2559 62 2625 572
rect 2751 62 2817 572
rect 2943 62 3009 572
rect 3135 62 3201 572
rect 3327 62 3393 572
rect 3519 62 3585 572
rect 3711 62 3777 572
rect 3903 62 3969 572
rect 4095 62 4161 572
rect 4287 62 4353 572
rect 4479 62 4545 572
rect 4671 62 4737 572
rect 4863 62 4929 572
rect 5055 62 5121 572
rect 5247 62 5313 572
rect 5439 62 5505 572
rect 5631 62 5697 572
rect 5823 62 5889 572
rect 6015 62 6081 572
rect 6207 62 6273 572
rect 6399 62 6465 572
rect 6591 62 6657 572
rect 6783 62 6849 572
rect 6975 62 7041 572
rect 7167 62 7233 572
rect 7359 62 7425 572
rect 7551 62 7617 572
rect 7743 62 7809 572
rect 7935 62 8001 572
rect 8127 62 8193 572
rect 8319 62 8385 572
rect 8511 62 8577 572
rect 8703 62 8769 572
rect 8895 62 8961 572
rect 9087 62 9153 572
rect 9279 62 9345 572
rect 9471 62 9537 572
rect 9663 62 9729 572
rect 9855 62 9921 572
rect 10047 62 10113 572
rect 10239 62 10305 572
rect 10431 62 10497 572
<< metal3 >>
rect -10507 572 -10421 582
rect -10507 62 -10497 572
rect -10431 62 -10421 572
rect -10507 52 -10421 62
rect -10315 572 -10229 582
rect -10315 62 -10305 572
rect -10239 62 -10229 572
rect -10315 52 -10229 62
rect -10123 572 -10037 582
rect -10123 62 -10113 572
rect -10047 62 -10037 572
rect -10123 52 -10037 62
rect -9931 572 -9845 582
rect -9931 62 -9921 572
rect -9855 62 -9845 572
rect -9931 52 -9845 62
rect -9739 572 -9653 582
rect -9739 62 -9729 572
rect -9663 62 -9653 572
rect -9739 52 -9653 62
rect -9547 572 -9461 582
rect -9547 62 -9537 572
rect -9471 62 -9461 572
rect -9547 52 -9461 62
rect -9355 572 -9269 582
rect -9355 62 -9345 572
rect -9279 62 -9269 572
rect -9355 52 -9269 62
rect -9163 572 -9077 582
rect -9163 62 -9153 572
rect -9087 62 -9077 572
rect -9163 52 -9077 62
rect -8971 572 -8885 582
rect -8971 62 -8961 572
rect -8895 62 -8885 572
rect -8971 52 -8885 62
rect -8779 572 -8693 582
rect -8779 62 -8769 572
rect -8703 62 -8693 572
rect -8779 52 -8693 62
rect -8587 572 -8501 582
rect -8587 62 -8577 572
rect -8511 62 -8501 572
rect -8587 52 -8501 62
rect -8395 572 -8309 582
rect -8395 62 -8385 572
rect -8319 62 -8309 572
rect -8395 52 -8309 62
rect -8203 572 -8117 582
rect -8203 62 -8193 572
rect -8127 62 -8117 572
rect -8203 52 -8117 62
rect -8011 572 -7925 582
rect -8011 62 -8001 572
rect -7935 62 -7925 572
rect -8011 52 -7925 62
rect -7819 572 -7733 582
rect -7819 62 -7809 572
rect -7743 62 -7733 572
rect -7819 52 -7733 62
rect -7627 572 -7541 582
rect -7627 62 -7617 572
rect -7551 62 -7541 572
rect -7627 52 -7541 62
rect -7435 572 -7349 582
rect -7435 62 -7425 572
rect -7359 62 -7349 572
rect -7435 52 -7349 62
rect -7243 572 -7157 582
rect -7243 62 -7233 572
rect -7167 62 -7157 572
rect -7243 52 -7157 62
rect -7051 572 -6965 582
rect -7051 62 -7041 572
rect -6975 62 -6965 572
rect -7051 52 -6965 62
rect -6859 572 -6773 582
rect -6859 62 -6849 572
rect -6783 62 -6773 572
rect -6859 52 -6773 62
rect -6667 572 -6581 582
rect -6667 62 -6657 572
rect -6591 62 -6581 572
rect -6667 52 -6581 62
rect -6475 572 -6389 582
rect -6475 62 -6465 572
rect -6399 62 -6389 572
rect -6475 52 -6389 62
rect -6283 572 -6197 582
rect -6283 62 -6273 572
rect -6207 62 -6197 572
rect -6283 52 -6197 62
rect -6091 572 -6005 582
rect -6091 62 -6081 572
rect -6015 62 -6005 572
rect -6091 52 -6005 62
rect -5899 572 -5813 582
rect -5899 62 -5889 572
rect -5823 62 -5813 572
rect -5899 52 -5813 62
rect -5707 572 -5621 582
rect -5707 62 -5697 572
rect -5631 62 -5621 572
rect -5707 52 -5621 62
rect -5515 572 -5429 582
rect -5515 62 -5505 572
rect -5439 62 -5429 572
rect -5515 52 -5429 62
rect -5323 572 -5237 582
rect -5323 62 -5313 572
rect -5247 62 -5237 572
rect -5323 52 -5237 62
rect -5131 572 -5045 582
rect -5131 62 -5121 572
rect -5055 62 -5045 572
rect -5131 52 -5045 62
rect -4939 572 -4853 582
rect -4939 62 -4929 572
rect -4863 62 -4853 572
rect -4939 52 -4853 62
rect -4747 572 -4661 582
rect -4747 62 -4737 572
rect -4671 62 -4661 572
rect -4747 52 -4661 62
rect -4555 572 -4469 582
rect -4555 62 -4545 572
rect -4479 62 -4469 572
rect -4555 52 -4469 62
rect -4363 572 -4277 582
rect -4363 62 -4353 572
rect -4287 62 -4277 572
rect -4363 52 -4277 62
rect -4171 572 -4085 582
rect -4171 62 -4161 572
rect -4095 62 -4085 572
rect -4171 52 -4085 62
rect -3979 572 -3893 582
rect -3979 62 -3969 572
rect -3903 62 -3893 572
rect -3979 52 -3893 62
rect -3787 572 -3701 582
rect -3787 62 -3777 572
rect -3711 62 -3701 572
rect -3787 52 -3701 62
rect -3595 572 -3509 582
rect -3595 62 -3585 572
rect -3519 62 -3509 572
rect -3595 52 -3509 62
rect -3403 572 -3317 582
rect -3403 62 -3393 572
rect -3327 62 -3317 572
rect -3403 52 -3317 62
rect -3211 572 -3125 582
rect -3211 62 -3201 572
rect -3135 62 -3125 572
rect -3211 52 -3125 62
rect -3019 572 -2933 582
rect -3019 62 -3009 572
rect -2943 62 -2933 572
rect -3019 52 -2933 62
rect -2827 572 -2741 582
rect -2827 62 -2817 572
rect -2751 62 -2741 572
rect -2827 52 -2741 62
rect -2635 572 -2549 582
rect -2635 62 -2625 572
rect -2559 62 -2549 572
rect -2635 52 -2549 62
rect -2443 572 -2357 582
rect -2443 62 -2433 572
rect -2367 62 -2357 572
rect -2443 52 -2357 62
rect -2251 572 -2165 582
rect -2251 62 -2241 572
rect -2175 62 -2165 572
rect -2251 52 -2165 62
rect -2059 572 -1973 582
rect -2059 62 -2049 572
rect -1983 62 -1973 572
rect -2059 52 -1973 62
rect -1867 572 -1781 582
rect -1867 62 -1857 572
rect -1791 62 -1781 572
rect -1867 52 -1781 62
rect -1675 572 -1589 582
rect -1675 62 -1665 572
rect -1599 62 -1589 572
rect -1675 52 -1589 62
rect -1483 572 -1397 582
rect -1483 62 -1473 572
rect -1407 62 -1397 572
rect -1483 52 -1397 62
rect -1291 572 -1205 582
rect -1291 62 -1281 572
rect -1215 62 -1205 572
rect -1291 52 -1205 62
rect -1099 572 -1013 582
rect -1099 62 -1089 572
rect -1023 62 -1013 572
rect -1099 52 -1013 62
rect -907 572 -821 582
rect -907 62 -897 572
rect -831 62 -821 572
rect -907 52 -821 62
rect -715 572 -629 582
rect -715 62 -705 572
rect -639 62 -629 572
rect -715 52 -629 62
rect -523 572 -437 582
rect -523 62 -513 572
rect -447 62 -437 572
rect -523 52 -437 62
rect -331 572 -245 582
rect -331 62 -321 572
rect -255 62 -245 572
rect -331 52 -245 62
rect -139 572 -53 582
rect -139 62 -129 572
rect -63 62 -53 572
rect -139 52 -53 62
rect 53 572 139 582
rect 53 62 63 572
rect 129 62 139 572
rect 53 52 139 62
rect 245 572 331 582
rect 245 62 255 572
rect 321 62 331 572
rect 245 52 331 62
rect 437 572 523 582
rect 437 62 447 572
rect 513 62 523 572
rect 437 52 523 62
rect 629 572 715 582
rect 629 62 639 572
rect 705 62 715 572
rect 629 52 715 62
rect 821 572 907 582
rect 821 62 831 572
rect 897 62 907 572
rect 821 52 907 62
rect 1013 572 1099 582
rect 1013 62 1023 572
rect 1089 62 1099 572
rect 1013 52 1099 62
rect 1205 572 1291 582
rect 1205 62 1215 572
rect 1281 62 1291 572
rect 1205 52 1291 62
rect 1397 572 1483 582
rect 1397 62 1407 572
rect 1473 62 1483 572
rect 1397 52 1483 62
rect 1589 572 1675 582
rect 1589 62 1599 572
rect 1665 62 1675 572
rect 1589 52 1675 62
rect 1781 572 1867 582
rect 1781 62 1791 572
rect 1857 62 1867 572
rect 1781 52 1867 62
rect 1973 572 2059 582
rect 1973 62 1983 572
rect 2049 62 2059 572
rect 1973 52 2059 62
rect 2165 572 2251 582
rect 2165 62 2175 572
rect 2241 62 2251 572
rect 2165 52 2251 62
rect 2357 572 2443 582
rect 2357 62 2367 572
rect 2433 62 2443 572
rect 2357 52 2443 62
rect 2549 572 2635 582
rect 2549 62 2559 572
rect 2625 62 2635 572
rect 2549 52 2635 62
rect 2741 572 2827 582
rect 2741 62 2751 572
rect 2817 62 2827 572
rect 2741 52 2827 62
rect 2933 572 3019 582
rect 2933 62 2943 572
rect 3009 62 3019 572
rect 2933 52 3019 62
rect 3125 572 3211 582
rect 3125 62 3135 572
rect 3201 62 3211 572
rect 3125 52 3211 62
rect 3317 572 3403 582
rect 3317 62 3327 572
rect 3393 62 3403 572
rect 3317 52 3403 62
rect 3509 572 3595 582
rect 3509 62 3519 572
rect 3585 62 3595 572
rect 3509 52 3595 62
rect 3701 572 3787 582
rect 3701 62 3711 572
rect 3777 62 3787 572
rect 3701 52 3787 62
rect 3893 572 3979 582
rect 3893 62 3903 572
rect 3969 62 3979 572
rect 3893 52 3979 62
rect 4085 572 4171 582
rect 4085 62 4095 572
rect 4161 62 4171 572
rect 4085 52 4171 62
rect 4277 572 4363 582
rect 4277 62 4287 572
rect 4353 62 4363 572
rect 4277 52 4363 62
rect 4469 572 4555 582
rect 4469 62 4479 572
rect 4545 62 4555 572
rect 4469 52 4555 62
rect 4661 572 4747 582
rect 4661 62 4671 572
rect 4737 62 4747 572
rect 4661 52 4747 62
rect 4853 572 4939 582
rect 4853 62 4863 572
rect 4929 62 4939 572
rect 4853 52 4939 62
rect 5045 572 5131 582
rect 5045 62 5055 572
rect 5121 62 5131 572
rect 5045 52 5131 62
rect 5237 572 5323 582
rect 5237 62 5247 572
rect 5313 62 5323 572
rect 5237 52 5323 62
rect 5429 572 5515 582
rect 5429 62 5439 572
rect 5505 62 5515 572
rect 5429 52 5515 62
rect 5621 572 5707 582
rect 5621 62 5631 572
rect 5697 62 5707 572
rect 5621 52 5707 62
rect 5813 572 5899 582
rect 5813 62 5823 572
rect 5889 62 5899 572
rect 5813 52 5899 62
rect 6005 572 6091 582
rect 6005 62 6015 572
rect 6081 62 6091 572
rect 6005 52 6091 62
rect 6197 572 6283 582
rect 6197 62 6207 572
rect 6273 62 6283 572
rect 6197 52 6283 62
rect 6389 572 6475 582
rect 6389 62 6399 572
rect 6465 62 6475 572
rect 6389 52 6475 62
rect 6581 572 6667 582
rect 6581 62 6591 572
rect 6657 62 6667 572
rect 6581 52 6667 62
rect 6773 572 6859 582
rect 6773 62 6783 572
rect 6849 62 6859 572
rect 6773 52 6859 62
rect 6965 572 7051 582
rect 6965 62 6975 572
rect 7041 62 7051 572
rect 6965 52 7051 62
rect 7157 572 7243 582
rect 7157 62 7167 572
rect 7233 62 7243 572
rect 7157 52 7243 62
rect 7349 572 7435 582
rect 7349 62 7359 572
rect 7425 62 7435 572
rect 7349 52 7435 62
rect 7541 572 7627 582
rect 7541 62 7551 572
rect 7617 62 7627 572
rect 7541 52 7627 62
rect 7733 572 7819 582
rect 7733 62 7743 572
rect 7809 62 7819 572
rect 7733 52 7819 62
rect 7925 572 8011 582
rect 7925 62 7935 572
rect 8001 62 8011 572
rect 7925 52 8011 62
rect 8117 572 8203 582
rect 8117 62 8127 572
rect 8193 62 8203 572
rect 8117 52 8203 62
rect 8309 572 8395 582
rect 8309 62 8319 572
rect 8385 62 8395 572
rect 8309 52 8395 62
rect 8501 572 8587 582
rect 8501 62 8511 572
rect 8577 62 8587 572
rect 8501 52 8587 62
rect 8693 572 8779 582
rect 8693 62 8703 572
rect 8769 62 8779 572
rect 8693 52 8779 62
rect 8885 572 8971 582
rect 8885 62 8895 572
rect 8961 62 8971 572
rect 8885 52 8971 62
rect 9077 572 9163 582
rect 9077 62 9087 572
rect 9153 62 9163 572
rect 9077 52 9163 62
rect 9269 572 9355 582
rect 9269 62 9279 572
rect 9345 62 9355 572
rect 9269 52 9355 62
rect 9461 572 9547 582
rect 9461 62 9471 572
rect 9537 62 9547 572
rect 9461 52 9547 62
rect 9653 572 9739 582
rect 9653 62 9663 572
rect 9729 62 9739 572
rect 9653 52 9739 62
rect 9845 572 9931 582
rect 9845 62 9855 572
rect 9921 62 9931 572
rect 9845 52 9931 62
rect 10037 572 10123 582
rect 10037 62 10047 572
rect 10113 62 10123 572
rect 10037 52 10123 62
rect 10229 572 10315 582
rect 10229 62 10239 572
rect 10305 62 10315 572
rect 10229 52 10315 62
rect 10421 572 10507 582
rect 10421 62 10431 572
rect 10497 62 10507 572
rect 10421 52 10507 62
<< via3 >>
rect -10497 62 -10431 572
rect -10305 62 -10239 572
rect -10113 62 -10047 572
rect -9921 62 -9855 572
rect -9729 62 -9663 572
rect -9537 62 -9471 572
rect -9345 62 -9279 572
rect -9153 62 -9087 572
rect -8961 62 -8895 572
rect -8769 62 -8703 572
rect -8577 62 -8511 572
rect -8385 62 -8319 572
rect -8193 62 -8127 572
rect -8001 62 -7935 572
rect -7809 62 -7743 572
rect -7617 62 -7551 572
rect -7425 62 -7359 572
rect -7233 62 -7167 572
rect -7041 62 -6975 572
rect -6849 62 -6783 572
rect -6657 62 -6591 572
rect -6465 62 -6399 572
rect -6273 62 -6207 572
rect -6081 62 -6015 572
rect -5889 62 -5823 572
rect -5697 62 -5631 572
rect -5505 62 -5439 572
rect -5313 62 -5247 572
rect -5121 62 -5055 572
rect -4929 62 -4863 572
rect -4737 62 -4671 572
rect -4545 62 -4479 572
rect -4353 62 -4287 572
rect -4161 62 -4095 572
rect -3969 62 -3903 572
rect -3777 62 -3711 572
rect -3585 62 -3519 572
rect -3393 62 -3327 572
rect -3201 62 -3135 572
rect -3009 62 -2943 572
rect -2817 62 -2751 572
rect -2625 62 -2559 572
rect -2433 62 -2367 572
rect -2241 62 -2175 572
rect -2049 62 -1983 572
rect -1857 62 -1791 572
rect -1665 62 -1599 572
rect -1473 62 -1407 572
rect -1281 62 -1215 572
rect -1089 62 -1023 572
rect -897 62 -831 572
rect -705 62 -639 572
rect -513 62 -447 572
rect -321 62 -255 572
rect -129 62 -63 572
rect 63 62 129 572
rect 255 62 321 572
rect 447 62 513 572
rect 639 62 705 572
rect 831 62 897 572
rect 1023 62 1089 572
rect 1215 62 1281 572
rect 1407 62 1473 572
rect 1599 62 1665 572
rect 1791 62 1857 572
rect 1983 62 2049 572
rect 2175 62 2241 572
rect 2367 62 2433 572
rect 2559 62 2625 572
rect 2751 62 2817 572
rect 2943 62 3009 572
rect 3135 62 3201 572
rect 3327 62 3393 572
rect 3519 62 3585 572
rect 3711 62 3777 572
rect 3903 62 3969 572
rect 4095 62 4161 572
rect 4287 62 4353 572
rect 4479 62 4545 572
rect 4671 62 4737 572
rect 4863 62 4929 572
rect 5055 62 5121 572
rect 5247 62 5313 572
rect 5439 62 5505 572
rect 5631 62 5697 572
rect 5823 62 5889 572
rect 6015 62 6081 572
rect 6207 62 6273 572
rect 6399 62 6465 572
rect 6591 62 6657 572
rect 6783 62 6849 572
rect 6975 62 7041 572
rect 7167 62 7233 572
rect 7359 62 7425 572
rect 7551 62 7617 572
rect 7743 62 7809 572
rect 7935 62 8001 572
rect 8127 62 8193 572
rect 8319 62 8385 572
rect 8511 62 8577 572
rect 8703 62 8769 572
rect 8895 62 8961 572
rect 9087 62 9153 572
rect 9279 62 9345 572
rect 9471 62 9537 572
rect 9663 62 9729 572
rect 9855 62 9921 572
rect 10047 62 10113 572
rect 10239 62 10305 572
rect 10431 62 10497 572
<< metal4 >>
rect -10507 572 -10421 582
rect -10507 62 -10497 572
rect -10431 62 -10421 572
rect -10507 52 -10421 62
rect -10315 572 -10229 582
rect -10315 62 -10305 572
rect -10239 62 -10229 572
rect -10315 52 -10229 62
rect -10123 572 -10037 582
rect -10123 62 -10113 572
rect -10047 62 -10037 572
rect -10123 52 -10037 62
rect -9931 572 -9845 582
rect -9931 62 -9921 572
rect -9855 62 -9845 572
rect -9931 52 -9845 62
rect -9739 572 -9653 582
rect -9739 62 -9729 572
rect -9663 62 -9653 572
rect -9739 52 -9653 62
rect -9547 572 -9461 582
rect -9547 62 -9537 572
rect -9471 62 -9461 572
rect -9547 52 -9461 62
rect -9355 572 -9269 582
rect -9355 62 -9345 572
rect -9279 62 -9269 572
rect -9355 52 -9269 62
rect -9163 572 -9077 582
rect -9163 62 -9153 572
rect -9087 62 -9077 572
rect -9163 52 -9077 62
rect -8971 572 -8885 582
rect -8971 62 -8961 572
rect -8895 62 -8885 572
rect -8971 52 -8885 62
rect -8779 572 -8693 582
rect -8779 62 -8769 572
rect -8703 62 -8693 572
rect -8779 52 -8693 62
rect -8587 572 -8501 582
rect -8587 62 -8577 572
rect -8511 62 -8501 572
rect -8587 52 -8501 62
rect -8395 572 -8309 582
rect -8395 62 -8385 572
rect -8319 62 -8309 572
rect -8395 52 -8309 62
rect -8203 572 -8117 582
rect -8203 62 -8193 572
rect -8127 62 -8117 572
rect -8203 52 -8117 62
rect -8011 572 -7925 582
rect -8011 62 -8001 572
rect -7935 62 -7925 572
rect -8011 52 -7925 62
rect -7819 572 -7733 582
rect -7819 62 -7809 572
rect -7743 62 -7733 572
rect -7819 52 -7733 62
rect -7627 572 -7541 582
rect -7627 62 -7617 572
rect -7551 62 -7541 572
rect -7627 52 -7541 62
rect -7435 572 -7349 582
rect -7435 62 -7425 572
rect -7359 62 -7349 572
rect -7435 52 -7349 62
rect -7243 572 -7157 582
rect -7243 62 -7233 572
rect -7167 62 -7157 572
rect -7243 52 -7157 62
rect -7051 572 -6965 582
rect -7051 62 -7041 572
rect -6975 62 -6965 572
rect -7051 52 -6965 62
rect -6859 572 -6773 582
rect -6859 62 -6849 572
rect -6783 62 -6773 572
rect -6859 52 -6773 62
rect -6667 572 -6581 582
rect -6667 62 -6657 572
rect -6591 62 -6581 572
rect -6667 52 -6581 62
rect -6475 572 -6389 582
rect -6475 62 -6465 572
rect -6399 62 -6389 572
rect -6475 52 -6389 62
rect -6283 572 -6197 582
rect -6283 62 -6273 572
rect -6207 62 -6197 572
rect -6283 52 -6197 62
rect -6091 572 -6005 582
rect -6091 62 -6081 572
rect -6015 62 -6005 572
rect -6091 52 -6005 62
rect -5899 572 -5813 582
rect -5899 62 -5889 572
rect -5823 62 -5813 572
rect -5899 52 -5813 62
rect -5707 572 -5621 582
rect -5707 62 -5697 572
rect -5631 62 -5621 572
rect -5707 52 -5621 62
rect -5515 572 -5429 582
rect -5515 62 -5505 572
rect -5439 62 -5429 572
rect -5515 52 -5429 62
rect -5323 572 -5237 582
rect -5323 62 -5313 572
rect -5247 62 -5237 572
rect -5323 52 -5237 62
rect -5131 572 -5045 582
rect -5131 62 -5121 572
rect -5055 62 -5045 572
rect -5131 52 -5045 62
rect -4939 572 -4853 582
rect -4939 62 -4929 572
rect -4863 62 -4853 572
rect -4939 52 -4853 62
rect -4747 572 -4661 582
rect -4747 62 -4737 572
rect -4671 62 -4661 572
rect -4747 52 -4661 62
rect -4555 572 -4469 582
rect -4555 62 -4545 572
rect -4479 62 -4469 572
rect -4555 52 -4469 62
rect -4363 572 -4277 582
rect -4363 62 -4353 572
rect -4287 62 -4277 572
rect -4363 52 -4277 62
rect -4171 572 -4085 582
rect -4171 62 -4161 572
rect -4095 62 -4085 572
rect -4171 52 -4085 62
rect -3979 572 -3893 582
rect -3979 62 -3969 572
rect -3903 62 -3893 572
rect -3979 52 -3893 62
rect -3787 572 -3701 582
rect -3787 62 -3777 572
rect -3711 62 -3701 572
rect -3787 52 -3701 62
rect -3595 572 -3509 582
rect -3595 62 -3585 572
rect -3519 62 -3509 572
rect -3595 52 -3509 62
rect -3403 572 -3317 582
rect -3403 62 -3393 572
rect -3327 62 -3317 572
rect -3403 52 -3317 62
rect -3211 572 -3125 582
rect -3211 62 -3201 572
rect -3135 62 -3125 572
rect -3211 52 -3125 62
rect -3019 572 -2933 582
rect -3019 62 -3009 572
rect -2943 62 -2933 572
rect -3019 52 -2933 62
rect -2827 572 -2741 582
rect -2827 62 -2817 572
rect -2751 62 -2741 572
rect -2827 52 -2741 62
rect -2635 572 -2549 582
rect -2635 62 -2625 572
rect -2559 62 -2549 572
rect -2635 52 -2549 62
rect -2443 572 -2357 582
rect -2443 62 -2433 572
rect -2367 62 -2357 572
rect -2443 52 -2357 62
rect -2251 572 -2165 582
rect -2251 62 -2241 572
rect -2175 62 -2165 572
rect -2251 52 -2165 62
rect -2059 572 -1973 582
rect -2059 62 -2049 572
rect -1983 62 -1973 572
rect -2059 52 -1973 62
rect -1867 572 -1781 582
rect -1867 62 -1857 572
rect -1791 62 -1781 572
rect -1867 52 -1781 62
rect -1675 572 -1589 582
rect -1675 62 -1665 572
rect -1599 62 -1589 572
rect -1675 52 -1589 62
rect -1483 572 -1397 582
rect -1483 62 -1473 572
rect -1407 62 -1397 572
rect -1483 52 -1397 62
rect -1291 572 -1205 582
rect -1291 62 -1281 572
rect -1215 62 -1205 572
rect -1291 52 -1205 62
rect -1099 572 -1013 582
rect -1099 62 -1089 572
rect -1023 62 -1013 572
rect -1099 52 -1013 62
rect -907 572 -821 582
rect -907 62 -897 572
rect -831 62 -821 572
rect -907 52 -821 62
rect -715 572 -629 582
rect -715 62 -705 572
rect -639 62 -629 572
rect -715 52 -629 62
rect -523 572 -437 582
rect -523 62 -513 572
rect -447 62 -437 572
rect -523 52 -437 62
rect -331 572 -245 582
rect -331 62 -321 572
rect -255 62 -245 572
rect -331 52 -245 62
rect -139 572 -53 582
rect -139 62 -129 572
rect -63 62 -53 572
rect -139 52 -53 62
rect 53 572 139 582
rect 53 62 63 572
rect 129 62 139 572
rect 53 52 139 62
rect 245 572 331 582
rect 245 62 255 572
rect 321 62 331 572
rect 245 52 331 62
rect 437 572 523 582
rect 437 62 447 572
rect 513 62 523 572
rect 437 52 523 62
rect 629 572 715 582
rect 629 62 639 572
rect 705 62 715 572
rect 629 52 715 62
rect 821 572 907 582
rect 821 62 831 572
rect 897 62 907 572
rect 821 52 907 62
rect 1013 572 1099 582
rect 1013 62 1023 572
rect 1089 62 1099 572
rect 1013 52 1099 62
rect 1205 572 1291 582
rect 1205 62 1215 572
rect 1281 62 1291 572
rect 1205 52 1291 62
rect 1397 572 1483 582
rect 1397 62 1407 572
rect 1473 62 1483 572
rect 1397 52 1483 62
rect 1589 572 1675 582
rect 1589 62 1599 572
rect 1665 62 1675 572
rect 1589 52 1675 62
rect 1781 572 1867 582
rect 1781 62 1791 572
rect 1857 62 1867 572
rect 1781 52 1867 62
rect 1973 572 2059 582
rect 1973 62 1983 572
rect 2049 62 2059 572
rect 1973 52 2059 62
rect 2165 572 2251 582
rect 2165 62 2175 572
rect 2241 62 2251 572
rect 2165 52 2251 62
rect 2357 572 2443 582
rect 2357 62 2367 572
rect 2433 62 2443 572
rect 2357 52 2443 62
rect 2549 572 2635 582
rect 2549 62 2559 572
rect 2625 62 2635 572
rect 2549 52 2635 62
rect 2741 572 2827 582
rect 2741 62 2751 572
rect 2817 62 2827 572
rect 2741 52 2827 62
rect 2933 572 3019 582
rect 2933 62 2943 572
rect 3009 62 3019 572
rect 2933 52 3019 62
rect 3125 572 3211 582
rect 3125 62 3135 572
rect 3201 62 3211 572
rect 3125 52 3211 62
rect 3317 572 3403 582
rect 3317 62 3327 572
rect 3393 62 3403 572
rect 3317 52 3403 62
rect 3509 572 3595 582
rect 3509 62 3519 572
rect 3585 62 3595 572
rect 3509 52 3595 62
rect 3701 572 3787 582
rect 3701 62 3711 572
rect 3777 62 3787 572
rect 3701 52 3787 62
rect 3893 572 3979 582
rect 3893 62 3903 572
rect 3969 62 3979 572
rect 3893 52 3979 62
rect 4085 572 4171 582
rect 4085 62 4095 572
rect 4161 62 4171 572
rect 4085 52 4171 62
rect 4277 572 4363 582
rect 4277 62 4287 572
rect 4353 62 4363 572
rect 4277 52 4363 62
rect 4469 572 4555 582
rect 4469 62 4479 572
rect 4545 62 4555 572
rect 4469 52 4555 62
rect 4661 572 4747 582
rect 4661 62 4671 572
rect 4737 62 4747 572
rect 4661 52 4747 62
rect 4853 572 4939 582
rect 4853 62 4863 572
rect 4929 62 4939 572
rect 4853 52 4939 62
rect 5045 572 5131 582
rect 5045 62 5055 572
rect 5121 62 5131 572
rect 5045 52 5131 62
rect 5237 572 5323 582
rect 5237 62 5247 572
rect 5313 62 5323 572
rect 5237 52 5323 62
rect 5429 572 5515 582
rect 5429 62 5439 572
rect 5505 62 5515 572
rect 5429 52 5515 62
rect 5621 572 5707 582
rect 5621 62 5631 572
rect 5697 62 5707 572
rect 5621 52 5707 62
rect 5813 572 5899 582
rect 5813 62 5823 572
rect 5889 62 5899 572
rect 5813 52 5899 62
rect 6005 572 6091 582
rect 6005 62 6015 572
rect 6081 62 6091 572
rect 6005 52 6091 62
rect 6197 572 6283 582
rect 6197 62 6207 572
rect 6273 62 6283 572
rect 6197 52 6283 62
rect 6389 572 6475 582
rect 6389 62 6399 572
rect 6465 62 6475 572
rect 6389 52 6475 62
rect 6581 572 6667 582
rect 6581 62 6591 572
rect 6657 62 6667 572
rect 6581 52 6667 62
rect 6773 572 6859 582
rect 6773 62 6783 572
rect 6849 62 6859 572
rect 6773 52 6859 62
rect 6965 572 7051 582
rect 6965 62 6975 572
rect 7041 62 7051 572
rect 6965 52 7051 62
rect 7157 572 7243 582
rect 7157 62 7167 572
rect 7233 62 7243 572
rect 7157 52 7243 62
rect 7349 572 7435 582
rect 7349 62 7359 572
rect 7425 62 7435 572
rect 7349 52 7435 62
rect 7541 572 7627 582
rect 7541 62 7551 572
rect 7617 62 7627 572
rect 7541 52 7627 62
rect 7733 572 7819 582
rect 7733 62 7743 572
rect 7809 62 7819 572
rect 7733 52 7819 62
rect 7925 572 8011 582
rect 7925 62 7935 572
rect 8001 62 8011 572
rect 7925 52 8011 62
rect 8117 572 8203 582
rect 8117 62 8127 572
rect 8193 62 8203 572
rect 8117 52 8203 62
rect 8309 572 8395 582
rect 8309 62 8319 572
rect 8385 62 8395 572
rect 8309 52 8395 62
rect 8501 572 8587 582
rect 8501 62 8511 572
rect 8577 62 8587 572
rect 8501 52 8587 62
rect 8693 572 8779 582
rect 8693 62 8703 572
rect 8769 62 8779 572
rect 8693 52 8779 62
rect 8885 572 8971 582
rect 8885 62 8895 572
rect 8961 62 8971 572
rect 8885 52 8971 62
rect 9077 572 9163 582
rect 9077 62 9087 572
rect 9153 62 9163 572
rect 9077 52 9163 62
rect 9269 572 9355 582
rect 9269 62 9279 572
rect 9345 62 9355 572
rect 9269 52 9355 62
rect 9461 572 9547 582
rect 9461 62 9471 572
rect 9537 62 9547 572
rect 9461 52 9547 62
rect 9653 572 9739 582
rect 9653 62 9663 572
rect 9729 62 9739 572
rect 9653 52 9739 62
rect 9845 572 9931 582
rect 9845 62 9855 572
rect 9921 62 9931 572
rect 9845 52 9931 62
rect 10037 572 10123 582
rect 10037 62 10047 572
rect 10113 62 10123 572
rect 10037 52 10123 62
rect 10229 572 10315 582
rect 10229 62 10239 572
rect 10305 62 10315 572
rect 10229 52 10315 62
rect 10421 572 10507 582
rect 10421 62 10431 572
rect 10497 62 10507 572
rect 10421 52 10507 62
<< properties >>
string FIXED_BBOX -10674 -866 10674 866
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 7 l 0.15 m 1 nf 220 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
