magic
tech sky130A
timestamp 1685741491
<< error_p >>
rect -2822 441 -2793 444
rect -2726 441 -2697 444
rect -2630 441 -2601 444
rect -2534 441 -2505 444
rect -2438 441 -2409 444
rect -2342 441 -2313 444
rect -2246 441 -2217 444
rect -2150 441 -2121 444
rect -2054 441 -2025 444
rect -1958 441 -1929 444
rect -1862 441 -1833 444
rect -1766 441 -1737 444
rect -1670 441 -1641 444
rect -1574 441 -1545 444
rect -1478 441 -1449 444
rect -1382 441 -1353 444
rect -1286 441 -1257 444
rect -1190 441 -1161 444
rect -1094 441 -1065 444
rect -998 441 -969 444
rect -902 441 -873 444
rect -806 441 -777 444
rect -710 441 -681 444
rect -614 441 -585 444
rect -518 441 -489 444
rect -422 441 -393 444
rect -326 441 -297 444
rect -230 441 -201 444
rect -134 441 -105 444
rect -38 441 -9 444
rect 57 441 86 444
rect 153 441 182 444
rect 249 441 278 444
rect 345 441 374 444
rect 441 441 470 444
rect 537 441 566 444
rect 633 441 662 444
rect 729 441 758 444
rect 825 441 854 444
rect 921 441 950 444
rect 1017 441 1046 444
rect 1113 441 1142 444
rect 1209 441 1238 444
rect 1305 441 1334 444
rect 1401 441 1430 444
rect 1497 441 1526 444
rect 1593 441 1622 444
rect 1689 441 1718 444
rect 1785 441 1814 444
rect 1881 441 1910 444
rect 1977 441 2006 444
rect 2073 441 2102 444
rect 2169 441 2198 444
rect 2265 441 2294 444
rect 2361 441 2390 444
rect 2457 441 2486 444
rect 2553 441 2582 444
rect 2649 441 2678 444
rect 2745 441 2774 444
rect 2841 441 2870 444
rect -2822 424 -2816 441
rect -2726 424 -2720 441
rect -2630 424 -2624 441
rect -2534 424 -2528 441
rect -2438 424 -2432 441
rect -2342 424 -2336 441
rect -2246 424 -2240 441
rect -2150 424 -2144 441
rect -2054 424 -2048 441
rect -1958 424 -1952 441
rect -1862 424 -1856 441
rect -1766 424 -1760 441
rect -1670 424 -1664 441
rect -1574 424 -1568 441
rect -1478 424 -1472 441
rect -1382 424 -1376 441
rect -1286 424 -1280 441
rect -1190 424 -1184 441
rect -1094 424 -1088 441
rect -998 424 -992 441
rect -902 424 -896 441
rect -806 424 -800 441
rect -710 424 -704 441
rect -614 424 -608 441
rect -518 424 -512 441
rect -422 424 -416 441
rect -326 424 -320 441
rect -230 424 -224 441
rect -134 424 -128 441
rect -38 424 -32 441
rect 57 424 63 441
rect 153 424 159 441
rect 249 424 255 441
rect 345 424 351 441
rect 441 424 447 441
rect 537 424 543 441
rect 633 424 639 441
rect 729 424 735 441
rect 825 424 831 441
rect 921 424 927 441
rect 1017 424 1023 441
rect 1113 424 1119 441
rect 1209 424 1215 441
rect 1305 424 1311 441
rect 1401 424 1407 441
rect 1497 424 1503 441
rect 1593 424 1599 441
rect 1689 424 1695 441
rect 1785 424 1791 441
rect 1881 424 1887 441
rect 1977 424 1983 441
rect 2073 424 2079 441
rect 2169 424 2175 441
rect 2265 424 2271 441
rect 2361 424 2367 441
rect 2457 424 2463 441
rect 2553 424 2559 441
rect 2649 424 2655 441
rect 2745 424 2751 441
rect 2841 424 2847 441
rect -2822 421 -2793 424
rect -2726 421 -2697 424
rect -2630 421 -2601 424
rect -2534 421 -2505 424
rect -2438 421 -2409 424
rect -2342 421 -2313 424
rect -2246 421 -2217 424
rect -2150 421 -2121 424
rect -2054 421 -2025 424
rect -1958 421 -1929 424
rect -1862 421 -1833 424
rect -1766 421 -1737 424
rect -1670 421 -1641 424
rect -1574 421 -1545 424
rect -1478 421 -1449 424
rect -1382 421 -1353 424
rect -1286 421 -1257 424
rect -1190 421 -1161 424
rect -1094 421 -1065 424
rect -998 421 -969 424
rect -902 421 -873 424
rect -806 421 -777 424
rect -710 421 -681 424
rect -614 421 -585 424
rect -518 421 -489 424
rect -422 421 -393 424
rect -326 421 -297 424
rect -230 421 -201 424
rect -134 421 -105 424
rect -38 421 -9 424
rect 57 421 86 424
rect 153 421 182 424
rect 249 421 278 424
rect 345 421 374 424
rect 441 421 470 424
rect 537 421 566 424
rect 633 421 662 424
rect 729 421 758 424
rect 825 421 854 424
rect 921 421 950 424
rect 1017 421 1046 424
rect 1113 421 1142 424
rect 1209 421 1238 424
rect 1305 421 1334 424
rect 1401 421 1430 424
rect 1497 421 1526 424
rect 1593 421 1622 424
rect 1689 421 1718 424
rect 1785 421 1814 424
rect 1881 421 1910 424
rect 1977 421 2006 424
rect 2073 421 2102 424
rect 2169 421 2198 424
rect 2265 421 2294 424
rect 2361 421 2390 424
rect 2457 421 2486 424
rect 2553 421 2582 424
rect 2649 421 2678 424
rect 2745 421 2774 424
rect 2841 421 2870 424
rect -2870 -425 -2841 -422
rect -2774 -425 -2745 -422
rect -2678 -425 -2649 -422
rect -2582 -425 -2553 -422
rect -2486 -425 -2457 -422
rect -2390 -425 -2361 -422
rect -2294 -425 -2265 -422
rect -2198 -425 -2169 -422
rect -2102 -425 -2073 -422
rect -2006 -425 -1977 -422
rect -1910 -425 -1881 -422
rect -1814 -425 -1785 -422
rect -1718 -425 -1689 -422
rect -1622 -425 -1593 -422
rect -1526 -425 -1497 -422
rect -1430 -425 -1401 -422
rect -1334 -425 -1305 -422
rect -1238 -425 -1209 -422
rect -1142 -424 -1113 -421
rect -1046 -424 -1017 -421
rect -950 -424 -921 -421
rect -854 -424 -825 -421
rect -758 -424 -729 -421
rect -662 -424 -633 -421
rect -566 -424 -537 -421
rect -470 -424 -441 -421
rect -374 -424 -345 -421
rect -278 -424 -249 -421
rect -182 -424 -153 -421
rect -86 -424 -57 -421
rect 9 -424 38 -421
rect 105 -424 134 -421
rect 201 -424 230 -421
rect 297 -424 326 -421
rect 393 -424 422 -421
rect 489 -424 518 -421
rect 585 -424 614 -421
rect 681 -424 710 -421
rect 777 -424 806 -421
rect 873 -424 902 -421
rect 969 -424 998 -421
rect 1065 -424 1094 -421
rect 1161 -424 1190 -421
rect 1257 -424 1286 -421
rect 1353 -424 1382 -421
rect 1449 -424 1478 -421
rect 1545 -424 1574 -421
rect 1641 -424 1670 -421
rect 1737 -424 1766 -421
rect 1833 -424 1862 -421
rect 1929 -424 1958 -421
rect 2025 -424 2054 -421
rect 2121 -424 2150 -421
rect 2217 -424 2246 -421
rect 2313 -424 2342 -421
rect 2409 -424 2438 -421
rect 2505 -424 2534 -421
rect 2601 -424 2630 -421
rect 2697 -424 2726 -421
rect 2793 -424 2822 -421
rect -2870 -442 -2864 -425
rect -2774 -442 -2768 -425
rect -2678 -442 -2672 -425
rect -2582 -442 -2576 -425
rect -2486 -442 -2480 -425
rect -2390 -442 -2384 -425
rect -2294 -442 -2288 -425
rect -2198 -442 -2192 -425
rect -2102 -442 -2096 -425
rect -2006 -442 -2000 -425
rect -1910 -442 -1904 -425
rect -1814 -442 -1808 -425
rect -1718 -442 -1712 -425
rect -1622 -442 -1616 -425
rect -1526 -442 -1520 -425
rect -1430 -442 -1424 -425
rect -1334 -442 -1328 -425
rect -1238 -442 -1232 -425
rect -1142 -441 -1136 -424
rect -1046 -441 -1040 -424
rect -950 -441 -944 -424
rect -854 -441 -848 -424
rect -758 -441 -752 -424
rect -662 -441 -656 -424
rect -566 -441 -560 -424
rect -470 -441 -464 -424
rect -374 -441 -368 -424
rect -278 -441 -272 -424
rect -182 -441 -176 -424
rect -86 -441 -80 -424
rect 9 -441 15 -424
rect 105 -441 111 -424
rect 201 -441 207 -424
rect 297 -441 303 -424
rect 393 -441 399 -424
rect 489 -441 495 -424
rect 585 -441 591 -424
rect 681 -441 687 -424
rect 777 -441 783 -424
rect 873 -441 879 -424
rect 969 -441 975 -424
rect 1065 -441 1071 -424
rect 1161 -441 1167 -424
rect 1257 -441 1263 -424
rect 1353 -441 1359 -424
rect 1449 -441 1455 -424
rect 1545 -441 1551 -424
rect 1641 -441 1647 -424
rect 1737 -441 1743 -424
rect 1833 -441 1839 -424
rect 1929 -441 1935 -424
rect 2025 -441 2031 -424
rect 2121 -441 2127 -424
rect 2217 -441 2223 -424
rect 2313 -441 2319 -424
rect 2409 -441 2415 -424
rect 2505 -441 2511 -424
rect 2601 -441 2607 -424
rect 2697 -441 2703 -424
rect 2793 -441 2799 -424
rect -2870 -445 -2841 -442
rect -2774 -445 -2745 -442
rect -2678 -445 -2649 -442
rect -2582 -445 -2553 -442
rect -2486 -445 -2457 -442
rect -2390 -445 -2361 -442
rect -2294 -445 -2265 -442
rect -2198 -445 -2169 -442
rect -2102 -445 -2073 -442
rect -2006 -445 -1977 -442
rect -1910 -445 -1881 -442
rect -1814 -445 -1785 -442
rect -1718 -445 -1689 -442
rect -1622 -445 -1593 -442
rect -1526 -445 -1497 -442
rect -1430 -445 -1401 -442
rect -1334 -445 -1305 -442
rect -1238 -445 -1209 -442
rect -1142 -444 -1113 -441
rect -1046 -444 -1017 -441
rect -950 -444 -921 -441
rect -854 -444 -825 -441
rect -758 -444 -729 -441
rect -662 -444 -633 -441
rect -566 -444 -537 -441
rect -470 -444 -441 -441
rect -374 -444 -345 -441
rect -278 -444 -249 -441
rect -182 -444 -153 -441
rect -86 -444 -57 -441
rect 9 -444 38 -441
rect 105 -444 134 -441
rect 201 -444 230 -441
rect 297 -444 326 -441
rect 393 -444 422 -441
rect 489 -444 518 -441
rect 585 -444 614 -441
rect 681 -444 710 -441
rect 777 -444 806 -441
rect 873 -444 902 -441
rect 969 -444 998 -441
rect 1065 -444 1094 -441
rect 1161 -444 1190 -441
rect 1257 -444 1286 -441
rect 1353 -444 1382 -441
rect 1449 -444 1478 -441
rect 1545 -444 1574 -441
rect 1641 -444 1670 -441
rect 1737 -444 1766 -441
rect 1833 -444 1862 -441
rect 1929 -444 1958 -441
rect 2025 -444 2054 -441
rect 2121 -444 2150 -441
rect 2217 -444 2246 -441
rect 2313 -444 2342 -441
rect 2409 -444 2438 -441
rect 2505 -444 2534 -441
rect 2601 -444 2630 -441
rect 2697 -444 2726 -441
rect 2793 -444 2822 -441
<< nwell >>
rect -2963 -509 2963 509
<< pmos >>
rect -2863 -400 -2848 400
rect -2815 -400 -2800 400
rect -2767 -400 -2752 400
rect -2719 -400 -2704 400
rect -2671 -400 -2656 400
rect -2623 -400 -2608 400
rect -2575 -400 -2560 400
rect -2527 -400 -2512 400
rect -2479 -400 -2464 400
rect -2431 -400 -2416 400
rect -2383 -400 -2368 400
rect -2335 -400 -2320 400
rect -2287 -400 -2272 400
rect -2239 -400 -2224 400
rect -2191 -400 -2176 400
rect -2143 -400 -2128 400
rect -2095 -400 -2080 400
rect -2047 -400 -2032 400
rect -1999 -400 -1984 400
rect -1951 -400 -1936 400
rect -1903 -400 -1888 400
rect -1855 -400 -1840 400
rect -1807 -400 -1792 400
rect -1759 -400 -1744 400
rect -1711 -400 -1696 400
rect -1663 -400 -1648 400
rect -1615 -400 -1600 400
rect -1567 -400 -1552 400
rect -1519 -400 -1504 400
rect -1471 -400 -1456 400
rect -1423 -400 -1408 400
rect -1375 -400 -1360 400
rect -1327 -400 -1312 400
rect -1279 -400 -1264 400
rect -1231 -400 -1216 400
rect -1183 -400 -1168 400
rect -1135 -400 -1120 400
rect -1087 -400 -1072 400
rect -1039 -400 -1024 400
rect -991 -400 -976 400
rect -943 -400 -928 400
rect -895 -400 -880 400
rect -847 -400 -832 400
rect -799 -400 -784 400
rect -751 -400 -736 400
rect -703 -400 -688 400
rect -655 -400 -640 400
rect -607 -400 -592 400
rect -559 -400 -544 400
rect -511 -400 -496 400
rect -463 -400 -448 400
rect -415 -400 -400 400
rect -367 -400 -352 400
rect -319 -400 -304 400
rect -271 -400 -256 400
rect -223 -400 -208 400
rect -175 -400 -160 400
rect -127 -400 -112 400
rect -79 -400 -64 400
rect -31 -400 -16 400
rect 16 -400 31 400
rect 64 -400 79 400
rect 112 -400 127 400
rect 160 -400 175 400
rect 208 -400 223 400
rect 256 -400 271 400
rect 304 -400 319 400
rect 352 -400 367 400
rect 400 -400 415 400
rect 448 -400 463 400
rect 496 -400 511 400
rect 544 -400 559 400
rect 592 -400 607 400
rect 640 -400 655 400
rect 688 -400 703 400
rect 736 -400 751 400
rect 784 -400 799 400
rect 832 -400 847 400
rect 880 -400 895 400
rect 928 -400 943 400
rect 976 -400 991 400
rect 1024 -400 1039 400
rect 1072 -400 1087 400
rect 1120 -400 1135 400
rect 1168 -400 1183 400
rect 1216 -400 1231 400
rect 1264 -400 1279 400
rect 1312 -400 1327 400
rect 1360 -400 1375 400
rect 1408 -400 1423 400
rect 1456 -400 1471 400
rect 1504 -400 1519 400
rect 1552 -400 1567 400
rect 1600 -400 1615 400
rect 1648 -400 1663 400
rect 1696 -400 1711 400
rect 1744 -400 1759 400
rect 1792 -400 1807 400
rect 1840 -400 1855 400
rect 1888 -400 1903 400
rect 1936 -400 1951 400
rect 1984 -400 1999 400
rect 2032 -400 2047 400
rect 2080 -400 2095 400
rect 2128 -400 2143 400
rect 2176 -400 2191 400
rect 2224 -400 2239 400
rect 2272 -400 2287 400
rect 2320 -400 2335 400
rect 2368 -400 2383 400
rect 2416 -400 2431 400
rect 2464 -400 2479 400
rect 2512 -400 2527 400
rect 2560 -400 2575 400
rect 2608 -400 2623 400
rect 2656 -400 2671 400
rect 2704 -400 2719 400
rect 2752 -400 2767 400
rect 2800 -400 2815 400
rect 2848 -400 2863 400
<< pdiff >>
rect -2894 394 -2863 400
rect -2894 -394 -2888 394
rect -2871 -394 -2863 394
rect -2894 -400 -2863 -394
rect -2848 394 -2815 400
rect -2848 -394 -2840 394
rect -2823 -394 -2815 394
rect -2848 -400 -2815 -394
rect -2800 394 -2767 400
rect -2800 -394 -2792 394
rect -2775 -394 -2767 394
rect -2800 -400 -2767 -394
rect -2752 394 -2719 400
rect -2752 -394 -2744 394
rect -2727 -394 -2719 394
rect -2752 -400 -2719 -394
rect -2704 394 -2671 400
rect -2704 -394 -2696 394
rect -2679 -394 -2671 394
rect -2704 -400 -2671 -394
rect -2656 394 -2623 400
rect -2656 -394 -2648 394
rect -2631 -394 -2623 394
rect -2656 -400 -2623 -394
rect -2608 394 -2575 400
rect -2608 -394 -2600 394
rect -2583 -394 -2575 394
rect -2608 -400 -2575 -394
rect -2560 394 -2527 400
rect -2560 -394 -2552 394
rect -2535 -394 -2527 394
rect -2560 -400 -2527 -394
rect -2512 394 -2479 400
rect -2512 -394 -2504 394
rect -2487 -394 -2479 394
rect -2512 -400 -2479 -394
rect -2464 394 -2431 400
rect -2464 -394 -2456 394
rect -2439 -394 -2431 394
rect -2464 -400 -2431 -394
rect -2416 394 -2383 400
rect -2416 -394 -2408 394
rect -2391 -394 -2383 394
rect -2416 -400 -2383 -394
rect -2368 394 -2335 400
rect -2368 -394 -2360 394
rect -2343 -394 -2335 394
rect -2368 -400 -2335 -394
rect -2320 394 -2287 400
rect -2320 -394 -2312 394
rect -2295 -394 -2287 394
rect -2320 -400 -2287 -394
rect -2272 394 -2239 400
rect -2272 -394 -2264 394
rect -2247 -394 -2239 394
rect -2272 -400 -2239 -394
rect -2224 394 -2191 400
rect -2224 -394 -2216 394
rect -2199 -394 -2191 394
rect -2224 -400 -2191 -394
rect -2176 394 -2143 400
rect -2176 -394 -2168 394
rect -2151 -394 -2143 394
rect -2176 -400 -2143 -394
rect -2128 394 -2095 400
rect -2128 -394 -2120 394
rect -2103 -394 -2095 394
rect -2128 -400 -2095 -394
rect -2080 394 -2047 400
rect -2080 -394 -2072 394
rect -2055 -394 -2047 394
rect -2080 -400 -2047 -394
rect -2032 394 -1999 400
rect -2032 -394 -2024 394
rect -2007 -394 -1999 394
rect -2032 -400 -1999 -394
rect -1984 394 -1951 400
rect -1984 -394 -1976 394
rect -1959 -394 -1951 394
rect -1984 -400 -1951 -394
rect -1936 394 -1903 400
rect -1936 -394 -1928 394
rect -1911 -394 -1903 394
rect -1936 -400 -1903 -394
rect -1888 394 -1855 400
rect -1888 -394 -1880 394
rect -1863 -394 -1855 394
rect -1888 -400 -1855 -394
rect -1840 394 -1807 400
rect -1840 -394 -1832 394
rect -1815 -394 -1807 394
rect -1840 -400 -1807 -394
rect -1792 394 -1759 400
rect -1792 -394 -1784 394
rect -1767 -394 -1759 394
rect -1792 -400 -1759 -394
rect -1744 394 -1711 400
rect -1744 -394 -1736 394
rect -1719 -394 -1711 394
rect -1744 -400 -1711 -394
rect -1696 394 -1663 400
rect -1696 -394 -1688 394
rect -1671 -394 -1663 394
rect -1696 -400 -1663 -394
rect -1648 394 -1615 400
rect -1648 -394 -1640 394
rect -1623 -394 -1615 394
rect -1648 -400 -1615 -394
rect -1600 394 -1567 400
rect -1600 -394 -1592 394
rect -1575 -394 -1567 394
rect -1600 -400 -1567 -394
rect -1552 394 -1519 400
rect -1552 -394 -1544 394
rect -1527 -394 -1519 394
rect -1552 -400 -1519 -394
rect -1504 394 -1471 400
rect -1504 -394 -1496 394
rect -1479 -394 -1471 394
rect -1504 -400 -1471 -394
rect -1456 394 -1423 400
rect -1456 -394 -1448 394
rect -1431 -394 -1423 394
rect -1456 -400 -1423 -394
rect -1408 394 -1375 400
rect -1408 -394 -1400 394
rect -1383 -394 -1375 394
rect -1408 -400 -1375 -394
rect -1360 394 -1327 400
rect -1360 -394 -1352 394
rect -1335 -394 -1327 394
rect -1360 -400 -1327 -394
rect -1312 394 -1279 400
rect -1312 -394 -1304 394
rect -1287 -394 -1279 394
rect -1312 -400 -1279 -394
rect -1264 394 -1231 400
rect -1264 -394 -1256 394
rect -1239 -394 -1231 394
rect -1264 -400 -1231 -394
rect -1216 394 -1183 400
rect -1216 -394 -1208 394
rect -1191 -394 -1183 394
rect -1216 -400 -1183 -394
rect -1168 394 -1135 400
rect -1168 -394 -1160 394
rect -1143 -394 -1135 394
rect -1168 -400 -1135 -394
rect -1120 394 -1087 400
rect -1120 -394 -1112 394
rect -1095 -394 -1087 394
rect -1120 -400 -1087 -394
rect -1072 394 -1039 400
rect -1072 -394 -1064 394
rect -1047 -394 -1039 394
rect -1072 -400 -1039 -394
rect -1024 394 -991 400
rect -1024 -394 -1016 394
rect -999 -394 -991 394
rect -1024 -400 -991 -394
rect -976 394 -943 400
rect -976 -394 -968 394
rect -951 -394 -943 394
rect -976 -400 -943 -394
rect -928 394 -895 400
rect -928 -394 -920 394
rect -903 -394 -895 394
rect -928 -400 -895 -394
rect -880 394 -847 400
rect -880 -394 -872 394
rect -855 -394 -847 394
rect -880 -400 -847 -394
rect -832 394 -799 400
rect -832 -394 -824 394
rect -807 -394 -799 394
rect -832 -400 -799 -394
rect -784 394 -751 400
rect -784 -394 -776 394
rect -759 -394 -751 394
rect -784 -400 -751 -394
rect -736 394 -703 400
rect -736 -394 -728 394
rect -711 -394 -703 394
rect -736 -400 -703 -394
rect -688 394 -655 400
rect -688 -394 -680 394
rect -663 -394 -655 394
rect -688 -400 -655 -394
rect -640 394 -607 400
rect -640 -394 -632 394
rect -615 -394 -607 394
rect -640 -400 -607 -394
rect -592 394 -559 400
rect -592 -394 -584 394
rect -567 -394 -559 394
rect -592 -400 -559 -394
rect -544 394 -511 400
rect -544 -394 -536 394
rect -519 -394 -511 394
rect -544 -400 -511 -394
rect -496 394 -463 400
rect -496 -394 -488 394
rect -471 -394 -463 394
rect -496 -400 -463 -394
rect -448 394 -415 400
rect -448 -394 -440 394
rect -423 -394 -415 394
rect -448 -400 -415 -394
rect -400 394 -367 400
rect -400 -394 -392 394
rect -375 -394 -367 394
rect -400 -400 -367 -394
rect -352 394 -319 400
rect -352 -394 -344 394
rect -327 -394 -319 394
rect -352 -400 -319 -394
rect -304 394 -271 400
rect -304 -394 -296 394
rect -279 -394 -271 394
rect -304 -400 -271 -394
rect -256 394 -223 400
rect -256 -394 -248 394
rect -231 -394 -223 394
rect -256 -400 -223 -394
rect -208 394 -175 400
rect -208 -394 -200 394
rect -183 -394 -175 394
rect -208 -400 -175 -394
rect -160 394 -127 400
rect -160 -394 -152 394
rect -135 -394 -127 394
rect -160 -400 -127 -394
rect -112 394 -79 400
rect -112 -394 -104 394
rect -87 -394 -79 394
rect -112 -400 -79 -394
rect -64 394 -31 400
rect -64 -394 -56 394
rect -39 -394 -31 394
rect -64 -400 -31 -394
rect -16 394 16 400
rect -16 -394 -8 394
rect 9 -394 16 394
rect -16 -400 16 -394
rect 31 394 64 400
rect 31 -394 39 394
rect 56 -394 64 394
rect 31 -400 64 -394
rect 79 394 112 400
rect 79 -394 87 394
rect 104 -394 112 394
rect 79 -400 112 -394
rect 127 394 160 400
rect 127 -394 135 394
rect 152 -394 160 394
rect 127 -400 160 -394
rect 175 394 208 400
rect 175 -394 183 394
rect 200 -394 208 394
rect 175 -400 208 -394
rect 223 394 256 400
rect 223 -394 231 394
rect 248 -394 256 394
rect 223 -400 256 -394
rect 271 394 304 400
rect 271 -394 279 394
rect 296 -394 304 394
rect 271 -400 304 -394
rect 319 394 352 400
rect 319 -394 327 394
rect 344 -394 352 394
rect 319 -400 352 -394
rect 367 394 400 400
rect 367 -394 375 394
rect 392 -394 400 394
rect 367 -400 400 -394
rect 415 394 448 400
rect 415 -394 423 394
rect 440 -394 448 394
rect 415 -400 448 -394
rect 463 394 496 400
rect 463 -394 471 394
rect 488 -394 496 394
rect 463 -400 496 -394
rect 511 394 544 400
rect 511 -394 519 394
rect 536 -394 544 394
rect 511 -400 544 -394
rect 559 394 592 400
rect 559 -394 567 394
rect 584 -394 592 394
rect 559 -400 592 -394
rect 607 394 640 400
rect 607 -394 615 394
rect 632 -394 640 394
rect 607 -400 640 -394
rect 655 394 688 400
rect 655 -394 663 394
rect 680 -394 688 394
rect 655 -400 688 -394
rect 703 394 736 400
rect 703 -394 711 394
rect 728 -394 736 394
rect 703 -400 736 -394
rect 751 394 784 400
rect 751 -394 759 394
rect 776 -394 784 394
rect 751 -400 784 -394
rect 799 394 832 400
rect 799 -394 807 394
rect 824 -394 832 394
rect 799 -400 832 -394
rect 847 394 880 400
rect 847 -394 855 394
rect 872 -394 880 394
rect 847 -400 880 -394
rect 895 394 928 400
rect 895 -394 903 394
rect 920 -394 928 394
rect 895 -400 928 -394
rect 943 394 976 400
rect 943 -394 951 394
rect 968 -394 976 394
rect 943 -400 976 -394
rect 991 394 1024 400
rect 991 -394 999 394
rect 1016 -394 1024 394
rect 991 -400 1024 -394
rect 1039 394 1072 400
rect 1039 -394 1047 394
rect 1064 -394 1072 394
rect 1039 -400 1072 -394
rect 1087 394 1120 400
rect 1087 -394 1095 394
rect 1112 -394 1120 394
rect 1087 -400 1120 -394
rect 1135 394 1168 400
rect 1135 -394 1143 394
rect 1160 -394 1168 394
rect 1135 -400 1168 -394
rect 1183 394 1216 400
rect 1183 -394 1191 394
rect 1208 -394 1216 394
rect 1183 -400 1216 -394
rect 1231 394 1264 400
rect 1231 -394 1239 394
rect 1256 -394 1264 394
rect 1231 -400 1264 -394
rect 1279 394 1312 400
rect 1279 -394 1287 394
rect 1304 -394 1312 394
rect 1279 -400 1312 -394
rect 1327 394 1360 400
rect 1327 -394 1335 394
rect 1352 -394 1360 394
rect 1327 -400 1360 -394
rect 1375 394 1408 400
rect 1375 -394 1383 394
rect 1400 -394 1408 394
rect 1375 -400 1408 -394
rect 1423 394 1456 400
rect 1423 -394 1431 394
rect 1448 -394 1456 394
rect 1423 -400 1456 -394
rect 1471 394 1504 400
rect 1471 -394 1479 394
rect 1496 -394 1504 394
rect 1471 -400 1504 -394
rect 1519 394 1552 400
rect 1519 -394 1527 394
rect 1544 -394 1552 394
rect 1519 -400 1552 -394
rect 1567 394 1600 400
rect 1567 -394 1575 394
rect 1592 -394 1600 394
rect 1567 -400 1600 -394
rect 1615 394 1648 400
rect 1615 -394 1623 394
rect 1640 -394 1648 394
rect 1615 -400 1648 -394
rect 1663 394 1696 400
rect 1663 -394 1671 394
rect 1688 -394 1696 394
rect 1663 -400 1696 -394
rect 1711 394 1744 400
rect 1711 -394 1719 394
rect 1736 -394 1744 394
rect 1711 -400 1744 -394
rect 1759 394 1792 400
rect 1759 -394 1767 394
rect 1784 -394 1792 394
rect 1759 -400 1792 -394
rect 1807 394 1840 400
rect 1807 -394 1815 394
rect 1832 -394 1840 394
rect 1807 -400 1840 -394
rect 1855 394 1888 400
rect 1855 -394 1863 394
rect 1880 -394 1888 394
rect 1855 -400 1888 -394
rect 1903 394 1936 400
rect 1903 -394 1911 394
rect 1928 -394 1936 394
rect 1903 -400 1936 -394
rect 1951 394 1984 400
rect 1951 -394 1959 394
rect 1976 -394 1984 394
rect 1951 -400 1984 -394
rect 1999 394 2032 400
rect 1999 -394 2007 394
rect 2024 -394 2032 394
rect 1999 -400 2032 -394
rect 2047 394 2080 400
rect 2047 -394 2055 394
rect 2072 -394 2080 394
rect 2047 -400 2080 -394
rect 2095 394 2128 400
rect 2095 -394 2103 394
rect 2120 -394 2128 394
rect 2095 -400 2128 -394
rect 2143 394 2176 400
rect 2143 -394 2151 394
rect 2168 -394 2176 394
rect 2143 -400 2176 -394
rect 2191 394 2224 400
rect 2191 -394 2199 394
rect 2216 -394 2224 394
rect 2191 -400 2224 -394
rect 2239 394 2272 400
rect 2239 -394 2247 394
rect 2264 -394 2272 394
rect 2239 -400 2272 -394
rect 2287 394 2320 400
rect 2287 -394 2295 394
rect 2312 -394 2320 394
rect 2287 -400 2320 -394
rect 2335 394 2368 400
rect 2335 -394 2343 394
rect 2360 -394 2368 394
rect 2335 -400 2368 -394
rect 2383 394 2416 400
rect 2383 -394 2391 394
rect 2408 -394 2416 394
rect 2383 -400 2416 -394
rect 2431 394 2464 400
rect 2431 -394 2439 394
rect 2456 -394 2464 394
rect 2431 -400 2464 -394
rect 2479 394 2512 400
rect 2479 -394 2487 394
rect 2504 -394 2512 394
rect 2479 -400 2512 -394
rect 2527 394 2560 400
rect 2527 -394 2535 394
rect 2552 -394 2560 394
rect 2527 -400 2560 -394
rect 2575 394 2608 400
rect 2575 -394 2583 394
rect 2600 -394 2608 394
rect 2575 -400 2608 -394
rect 2623 394 2656 400
rect 2623 -394 2631 394
rect 2648 -394 2656 394
rect 2623 -400 2656 -394
rect 2671 394 2704 400
rect 2671 -394 2679 394
rect 2696 -394 2704 394
rect 2671 -400 2704 -394
rect 2719 394 2752 400
rect 2719 -394 2727 394
rect 2744 -394 2752 394
rect 2719 -400 2752 -394
rect 2767 394 2800 400
rect 2767 -394 2775 394
rect 2792 -394 2800 394
rect 2767 -400 2800 -394
rect 2815 394 2848 400
rect 2815 -394 2823 394
rect 2840 -394 2848 394
rect 2815 -400 2848 -394
rect 2863 394 2894 400
rect 2863 -394 2871 394
rect 2888 -394 2894 394
rect 2863 -400 2894 -394
<< pdiffc >>
rect -2888 -394 -2871 394
rect -2840 -394 -2823 394
rect -2792 -394 -2775 394
rect -2744 -394 -2727 394
rect -2696 -394 -2679 394
rect -2648 -394 -2631 394
rect -2600 -394 -2583 394
rect -2552 -394 -2535 394
rect -2504 -394 -2487 394
rect -2456 -394 -2439 394
rect -2408 -394 -2391 394
rect -2360 -394 -2343 394
rect -2312 -394 -2295 394
rect -2264 -394 -2247 394
rect -2216 -394 -2199 394
rect -2168 -394 -2151 394
rect -2120 -394 -2103 394
rect -2072 -394 -2055 394
rect -2024 -394 -2007 394
rect -1976 -394 -1959 394
rect -1928 -394 -1911 394
rect -1880 -394 -1863 394
rect -1832 -394 -1815 394
rect -1784 -394 -1767 394
rect -1736 -394 -1719 394
rect -1688 -394 -1671 394
rect -1640 -394 -1623 394
rect -1592 -394 -1575 394
rect -1544 -394 -1527 394
rect -1496 -394 -1479 394
rect -1448 -394 -1431 394
rect -1400 -394 -1383 394
rect -1352 -394 -1335 394
rect -1304 -394 -1287 394
rect -1256 -394 -1239 394
rect -1208 -394 -1191 394
rect -1160 -394 -1143 394
rect -1112 -394 -1095 394
rect -1064 -394 -1047 394
rect -1016 -394 -999 394
rect -968 -394 -951 394
rect -920 -394 -903 394
rect -872 -394 -855 394
rect -824 -394 -807 394
rect -776 -394 -759 394
rect -728 -394 -711 394
rect -680 -394 -663 394
rect -632 -394 -615 394
rect -584 -394 -567 394
rect -536 -394 -519 394
rect -488 -394 -471 394
rect -440 -394 -423 394
rect -392 -394 -375 394
rect -344 -394 -327 394
rect -296 -394 -279 394
rect -248 -394 -231 394
rect -200 -394 -183 394
rect -152 -394 -135 394
rect -104 -394 -87 394
rect -56 -394 -39 394
rect -8 -394 9 394
rect 39 -394 56 394
rect 87 -394 104 394
rect 135 -394 152 394
rect 183 -394 200 394
rect 231 -394 248 394
rect 279 -394 296 394
rect 327 -394 344 394
rect 375 -394 392 394
rect 423 -394 440 394
rect 471 -394 488 394
rect 519 -394 536 394
rect 567 -394 584 394
rect 615 -394 632 394
rect 663 -394 680 394
rect 711 -394 728 394
rect 759 -394 776 394
rect 807 -394 824 394
rect 855 -394 872 394
rect 903 -394 920 394
rect 951 -394 968 394
rect 999 -394 1016 394
rect 1047 -394 1064 394
rect 1095 -394 1112 394
rect 1143 -394 1160 394
rect 1191 -394 1208 394
rect 1239 -394 1256 394
rect 1287 -394 1304 394
rect 1335 -394 1352 394
rect 1383 -394 1400 394
rect 1431 -394 1448 394
rect 1479 -394 1496 394
rect 1527 -394 1544 394
rect 1575 -394 1592 394
rect 1623 -394 1640 394
rect 1671 -394 1688 394
rect 1719 -394 1736 394
rect 1767 -394 1784 394
rect 1815 -394 1832 394
rect 1863 -394 1880 394
rect 1911 -394 1928 394
rect 1959 -394 1976 394
rect 2007 -394 2024 394
rect 2055 -394 2072 394
rect 2103 -394 2120 394
rect 2151 -394 2168 394
rect 2199 -394 2216 394
rect 2247 -394 2264 394
rect 2295 -394 2312 394
rect 2343 -394 2360 394
rect 2391 -394 2408 394
rect 2439 -394 2456 394
rect 2487 -394 2504 394
rect 2535 -394 2552 394
rect 2583 -394 2600 394
rect 2631 -394 2648 394
rect 2679 -394 2696 394
rect 2727 -394 2744 394
rect 2775 -394 2792 394
rect 2823 -394 2840 394
rect 2871 -394 2888 394
<< nsubdiff >>
rect -2945 474 -2897 491
rect 2897 474 2945 491
rect -2945 443 -2928 474
rect 2928 443 2945 474
rect -2945 -474 -2928 -443
rect 2928 -474 2945 -443
rect -2945 -491 -2897 -474
rect 2897 -491 2945 -474
<< nsubdiffcont >>
rect -2897 474 2897 491
rect -2945 -443 -2928 443
rect 2928 -443 2945 443
rect -2897 -491 2897 -474
<< poly >>
rect -2824 441 -2791 449
rect -2824 424 -2816 441
rect -2799 424 -2791 441
rect -2824 416 -2791 424
rect -2728 441 -2695 449
rect -2728 424 -2720 441
rect -2703 424 -2695 441
rect -2728 416 -2695 424
rect -2632 441 -2599 449
rect -2632 424 -2624 441
rect -2607 424 -2599 441
rect -2632 416 -2599 424
rect -2536 441 -2503 449
rect -2536 424 -2528 441
rect -2511 424 -2503 441
rect -2536 416 -2503 424
rect -2440 441 -2407 449
rect -2440 424 -2432 441
rect -2415 424 -2407 441
rect -2440 416 -2407 424
rect -2344 441 -2311 449
rect -2344 424 -2336 441
rect -2319 424 -2311 441
rect -2344 416 -2311 424
rect -2248 441 -2215 449
rect -2248 424 -2240 441
rect -2223 424 -2215 441
rect -2248 416 -2215 424
rect -2152 441 -2119 449
rect -2152 424 -2144 441
rect -2127 424 -2119 441
rect -2152 416 -2119 424
rect -2056 441 -2023 449
rect -2056 424 -2048 441
rect -2031 424 -2023 441
rect -2056 416 -2023 424
rect -1960 441 -1927 449
rect -1960 424 -1952 441
rect -1935 424 -1927 441
rect -1960 416 -1927 424
rect -1864 441 -1831 449
rect -1864 424 -1856 441
rect -1839 424 -1831 441
rect -1864 416 -1831 424
rect -1768 441 -1735 449
rect -1768 424 -1760 441
rect -1743 424 -1735 441
rect -1768 416 -1735 424
rect -1672 441 -1639 449
rect -1672 424 -1664 441
rect -1647 424 -1639 441
rect -1672 416 -1639 424
rect -1576 441 -1543 449
rect -1576 424 -1568 441
rect -1551 424 -1543 441
rect -1576 416 -1543 424
rect -1480 441 -1447 449
rect -1480 424 -1472 441
rect -1455 424 -1447 441
rect -1480 416 -1447 424
rect -1384 441 -1351 449
rect -1384 424 -1376 441
rect -1359 424 -1351 441
rect -1384 416 -1351 424
rect -1288 441 -1255 449
rect -1288 424 -1280 441
rect -1263 424 -1255 441
rect -1288 416 -1255 424
rect -1192 441 -1159 449
rect -1192 424 -1184 441
rect -1167 424 -1159 441
rect -1192 416 -1159 424
rect -1096 441 -1063 449
rect -1096 424 -1088 441
rect -1071 424 -1063 441
rect -1096 416 -1063 424
rect -1000 441 -967 449
rect -1000 424 -992 441
rect -975 424 -967 441
rect -1000 416 -967 424
rect -904 441 -871 449
rect -904 424 -896 441
rect -879 424 -871 441
rect -904 416 -871 424
rect -808 441 -775 449
rect -808 424 -800 441
rect -783 424 -775 441
rect -808 416 -775 424
rect -712 441 -679 449
rect -712 424 -704 441
rect -687 424 -679 441
rect -712 416 -679 424
rect -616 441 -583 449
rect -616 424 -608 441
rect -591 424 -583 441
rect -616 416 -583 424
rect -520 441 -487 449
rect -520 424 -512 441
rect -495 424 -487 441
rect -520 416 -487 424
rect -424 441 -391 449
rect -424 424 -416 441
rect -399 424 -391 441
rect -424 416 -391 424
rect -328 441 -295 449
rect -328 424 -320 441
rect -303 424 -295 441
rect -328 416 -295 424
rect -232 441 -199 449
rect -232 424 -224 441
rect -207 424 -199 441
rect -232 416 -199 424
rect -136 441 -103 449
rect -136 424 -128 441
rect -111 424 -103 441
rect -136 416 -103 424
rect -40 441 -7 449
rect -40 424 -32 441
rect -15 424 -7 441
rect -40 416 -7 424
rect 55 441 88 449
rect 55 424 63 441
rect 80 424 88 441
rect 55 416 88 424
rect 151 441 184 449
rect 151 424 159 441
rect 176 424 184 441
rect 151 416 184 424
rect 247 441 280 449
rect 247 424 255 441
rect 272 424 280 441
rect 247 416 280 424
rect 343 441 376 449
rect 343 424 351 441
rect 368 424 376 441
rect 343 416 376 424
rect 439 441 472 449
rect 439 424 447 441
rect 464 424 472 441
rect 439 416 472 424
rect 535 441 568 449
rect 535 424 543 441
rect 560 424 568 441
rect 535 416 568 424
rect 631 441 664 449
rect 631 424 639 441
rect 656 424 664 441
rect 631 416 664 424
rect 727 441 760 449
rect 727 424 735 441
rect 752 424 760 441
rect 727 416 760 424
rect 823 441 856 449
rect 823 424 831 441
rect 848 424 856 441
rect 823 416 856 424
rect 919 441 952 449
rect 919 424 927 441
rect 944 424 952 441
rect 919 416 952 424
rect 1015 441 1048 449
rect 1015 424 1023 441
rect 1040 424 1048 441
rect 1015 416 1048 424
rect 1111 441 1144 449
rect 1111 424 1119 441
rect 1136 424 1144 441
rect 1111 416 1144 424
rect 1207 441 1240 449
rect 1207 424 1215 441
rect 1232 424 1240 441
rect 1207 416 1240 424
rect 1303 441 1336 449
rect 1303 424 1311 441
rect 1328 424 1336 441
rect 1303 416 1336 424
rect 1399 441 1432 449
rect 1399 424 1407 441
rect 1424 424 1432 441
rect 1399 416 1432 424
rect 1495 441 1528 449
rect 1495 424 1503 441
rect 1520 424 1528 441
rect 1495 416 1528 424
rect 1591 441 1624 449
rect 1591 424 1599 441
rect 1616 424 1624 441
rect 1591 416 1624 424
rect 1687 441 1720 449
rect 1687 424 1695 441
rect 1712 424 1720 441
rect 1687 416 1720 424
rect 1783 441 1816 449
rect 1783 424 1791 441
rect 1808 424 1816 441
rect 1783 416 1816 424
rect 1879 441 1912 449
rect 1879 424 1887 441
rect 1904 424 1912 441
rect 1879 416 1912 424
rect 1975 441 2008 449
rect 1975 424 1983 441
rect 2000 424 2008 441
rect 1975 416 2008 424
rect 2071 441 2104 449
rect 2071 424 2079 441
rect 2096 424 2104 441
rect 2071 416 2104 424
rect 2167 441 2200 449
rect 2167 424 2175 441
rect 2192 424 2200 441
rect 2167 416 2200 424
rect 2263 441 2296 449
rect 2263 424 2271 441
rect 2288 424 2296 441
rect 2263 416 2296 424
rect 2359 441 2392 449
rect 2359 424 2367 441
rect 2384 424 2392 441
rect 2359 416 2392 424
rect 2455 441 2488 449
rect 2455 424 2463 441
rect 2480 424 2488 441
rect 2455 416 2488 424
rect 2551 441 2584 449
rect 2551 424 2559 441
rect 2576 424 2584 441
rect 2551 416 2584 424
rect 2647 441 2680 449
rect 2647 424 2655 441
rect 2672 424 2680 441
rect 2647 416 2680 424
rect 2743 441 2776 449
rect 2743 424 2751 441
rect 2768 424 2776 441
rect 2743 416 2776 424
rect 2839 441 2872 449
rect 2839 424 2847 441
rect 2864 424 2872 441
rect 2839 416 2872 424
rect -2863 400 -2848 413
rect -2815 400 -2800 416
rect -2767 400 -2752 413
rect -2719 400 -2704 416
rect -2671 400 -2656 413
rect -2623 400 -2608 416
rect -2575 400 -2560 413
rect -2527 400 -2512 416
rect -2479 400 -2464 413
rect -2431 400 -2416 416
rect -2383 400 -2368 413
rect -2335 400 -2320 416
rect -2287 400 -2272 413
rect -2239 400 -2224 416
rect -2191 400 -2176 413
rect -2143 400 -2128 416
rect -2095 400 -2080 413
rect -2047 400 -2032 416
rect -1999 400 -1984 413
rect -1951 400 -1936 416
rect -1903 400 -1888 413
rect -1855 400 -1840 416
rect -1807 400 -1792 413
rect -1759 400 -1744 416
rect -1711 400 -1696 413
rect -1663 400 -1648 416
rect -1615 400 -1600 413
rect -1567 400 -1552 416
rect -1519 400 -1504 413
rect -1471 400 -1456 416
rect -1423 400 -1408 413
rect -1375 400 -1360 416
rect -1327 400 -1312 413
rect -1279 400 -1264 416
rect -1231 400 -1216 413
rect -1183 400 -1168 416
rect -1135 400 -1120 413
rect -1087 400 -1072 416
rect -1039 400 -1024 413
rect -991 400 -976 416
rect -943 400 -928 413
rect -895 400 -880 416
rect -847 400 -832 413
rect -799 400 -784 416
rect -751 400 -736 413
rect -703 400 -688 416
rect -655 400 -640 413
rect -607 400 -592 416
rect -559 400 -544 413
rect -511 400 -496 416
rect -463 400 -448 413
rect -415 400 -400 416
rect -367 400 -352 413
rect -319 400 -304 416
rect -271 400 -256 413
rect -223 400 -208 416
rect -175 400 -160 413
rect -127 400 -112 416
rect -79 400 -64 413
rect -31 400 -16 416
rect 16 400 31 413
rect 64 400 79 416
rect 112 400 127 413
rect 160 400 175 416
rect 208 400 223 413
rect 256 400 271 416
rect 304 400 319 413
rect 352 400 367 416
rect 400 400 415 413
rect 448 400 463 416
rect 496 400 511 413
rect 544 400 559 416
rect 592 400 607 413
rect 640 400 655 416
rect 688 400 703 413
rect 736 400 751 416
rect 784 400 799 413
rect 832 400 847 416
rect 880 400 895 413
rect 928 400 943 416
rect 976 400 991 413
rect 1024 400 1039 416
rect 1072 400 1087 413
rect 1120 400 1135 416
rect 1168 400 1183 413
rect 1216 400 1231 416
rect 1264 400 1279 413
rect 1312 400 1327 416
rect 1360 400 1375 413
rect 1408 400 1423 416
rect 1456 400 1471 413
rect 1504 400 1519 416
rect 1552 400 1567 413
rect 1600 400 1615 416
rect 1648 400 1663 413
rect 1696 400 1711 416
rect 1744 400 1759 413
rect 1792 400 1807 416
rect 1840 400 1855 413
rect 1888 400 1903 416
rect 1936 400 1951 413
rect 1984 400 1999 416
rect 2032 400 2047 413
rect 2080 400 2095 416
rect 2128 400 2143 413
rect 2176 400 2191 416
rect 2224 400 2239 413
rect 2272 400 2287 416
rect 2320 400 2335 413
rect 2368 400 2383 416
rect 2416 400 2431 413
rect 2464 400 2479 416
rect 2512 400 2527 413
rect 2560 400 2575 416
rect 2608 400 2623 413
rect 2656 400 2671 416
rect 2704 400 2719 413
rect 2752 400 2767 416
rect 2800 400 2815 413
rect 2848 400 2863 416
rect -2863 -417 -2848 -400
rect -2815 -413 -2800 -400
rect -2767 -417 -2752 -400
rect -2719 -413 -2704 -400
rect -2671 -417 -2656 -400
rect -2623 -413 -2608 -400
rect -2575 -417 -2560 -400
rect -2527 -413 -2512 -400
rect -2479 -417 -2464 -400
rect -2431 -413 -2416 -400
rect -2383 -417 -2368 -400
rect -2335 -413 -2320 -400
rect -2287 -417 -2272 -400
rect -2239 -413 -2224 -400
rect -2191 -417 -2176 -400
rect -2143 -413 -2128 -400
rect -2095 -417 -2080 -400
rect -2047 -413 -2032 -400
rect -1999 -417 -1984 -400
rect -1951 -413 -1936 -400
rect -1903 -417 -1888 -400
rect -1855 -413 -1840 -400
rect -1807 -417 -1792 -400
rect -1759 -413 -1744 -400
rect -1711 -417 -1696 -400
rect -1663 -413 -1648 -400
rect -1615 -417 -1600 -400
rect -1567 -413 -1552 -400
rect -1519 -417 -1504 -400
rect -1471 -413 -1456 -400
rect -1423 -417 -1408 -400
rect -1375 -413 -1360 -400
rect -1327 -417 -1312 -400
rect -1279 -413 -1264 -400
rect -1231 -417 -1216 -400
rect -1183 -413 -1168 -400
rect -1135 -416 -1120 -400
rect -1087 -413 -1072 -400
rect -1039 -416 -1024 -400
rect -991 -413 -976 -400
rect -943 -416 -928 -400
rect -895 -413 -880 -400
rect -847 -416 -832 -400
rect -799 -413 -784 -400
rect -751 -416 -736 -400
rect -703 -413 -688 -400
rect -655 -416 -640 -400
rect -607 -413 -592 -400
rect -559 -416 -544 -400
rect -511 -413 -496 -400
rect -463 -416 -448 -400
rect -415 -413 -400 -400
rect -367 -416 -352 -400
rect -319 -413 -304 -400
rect -271 -416 -256 -400
rect -223 -413 -208 -400
rect -175 -416 -160 -400
rect -127 -413 -112 -400
rect -79 -416 -64 -400
rect -31 -413 -16 -400
rect 16 -416 31 -400
rect 64 -413 79 -400
rect 112 -416 127 -400
rect 160 -413 175 -400
rect 208 -416 223 -400
rect 256 -413 271 -400
rect 304 -416 319 -400
rect 352 -413 367 -400
rect 400 -416 415 -400
rect 448 -413 463 -400
rect 496 -416 511 -400
rect 544 -413 559 -400
rect 592 -416 607 -400
rect 640 -413 655 -400
rect 688 -416 703 -400
rect 736 -413 751 -400
rect 784 -416 799 -400
rect 832 -413 847 -400
rect 880 -416 895 -400
rect 928 -413 943 -400
rect 976 -416 991 -400
rect 1024 -413 1039 -400
rect 1072 -416 1087 -400
rect 1120 -413 1135 -400
rect 1168 -416 1183 -400
rect 1216 -413 1231 -400
rect 1264 -416 1279 -400
rect 1312 -413 1327 -400
rect 1360 -416 1375 -400
rect 1408 -413 1423 -400
rect 1456 -416 1471 -400
rect 1504 -413 1519 -400
rect 1552 -416 1567 -400
rect 1600 -413 1615 -400
rect 1648 -416 1663 -400
rect 1696 -413 1711 -400
rect 1744 -416 1759 -400
rect 1792 -413 1807 -400
rect 1840 -416 1855 -400
rect 1888 -413 1903 -400
rect 1936 -416 1951 -400
rect 1984 -413 1999 -400
rect 2032 -416 2047 -400
rect 2080 -413 2095 -400
rect 2128 -416 2143 -400
rect 2176 -413 2191 -400
rect 2224 -416 2239 -400
rect 2272 -413 2287 -400
rect 2320 -416 2335 -400
rect 2368 -413 2383 -400
rect 2416 -416 2431 -400
rect 2464 -413 2479 -400
rect 2512 -416 2527 -400
rect 2560 -413 2575 -400
rect 2608 -416 2623 -400
rect 2656 -413 2671 -400
rect 2704 -416 2719 -400
rect 2752 -413 2767 -400
rect 2800 -416 2815 -400
rect 2848 -413 2863 -400
rect -2872 -425 -2839 -417
rect -2872 -442 -2864 -425
rect -2847 -442 -2839 -425
rect -2872 -450 -2839 -442
rect -2776 -425 -2743 -417
rect -2776 -442 -2768 -425
rect -2751 -442 -2743 -425
rect -2776 -450 -2743 -442
rect -2680 -425 -2647 -417
rect -2680 -442 -2672 -425
rect -2655 -442 -2647 -425
rect -2680 -450 -2647 -442
rect -2584 -425 -2551 -417
rect -2584 -442 -2576 -425
rect -2559 -442 -2551 -425
rect -2584 -450 -2551 -442
rect -2488 -425 -2455 -417
rect -2488 -442 -2480 -425
rect -2463 -442 -2455 -425
rect -2488 -450 -2455 -442
rect -2392 -425 -2359 -417
rect -2392 -442 -2384 -425
rect -2367 -442 -2359 -425
rect -2392 -450 -2359 -442
rect -2296 -425 -2263 -417
rect -2296 -442 -2288 -425
rect -2271 -442 -2263 -425
rect -2296 -450 -2263 -442
rect -2200 -425 -2167 -417
rect -2200 -442 -2192 -425
rect -2175 -442 -2167 -425
rect -2200 -450 -2167 -442
rect -2104 -425 -2071 -417
rect -2104 -442 -2096 -425
rect -2079 -442 -2071 -425
rect -2104 -450 -2071 -442
rect -2008 -425 -1975 -417
rect -2008 -442 -2000 -425
rect -1983 -442 -1975 -425
rect -2008 -450 -1975 -442
rect -1912 -425 -1879 -417
rect -1912 -442 -1904 -425
rect -1887 -442 -1879 -425
rect -1912 -450 -1879 -442
rect -1816 -425 -1783 -417
rect -1816 -442 -1808 -425
rect -1791 -442 -1783 -425
rect -1816 -450 -1783 -442
rect -1720 -425 -1687 -417
rect -1720 -442 -1712 -425
rect -1695 -442 -1687 -425
rect -1720 -450 -1687 -442
rect -1624 -425 -1591 -417
rect -1624 -442 -1616 -425
rect -1599 -442 -1591 -425
rect -1624 -450 -1591 -442
rect -1528 -425 -1495 -417
rect -1528 -442 -1520 -425
rect -1503 -442 -1495 -425
rect -1528 -450 -1495 -442
rect -1432 -425 -1399 -417
rect -1432 -442 -1424 -425
rect -1407 -442 -1399 -425
rect -1432 -450 -1399 -442
rect -1336 -425 -1303 -417
rect -1336 -442 -1328 -425
rect -1311 -442 -1303 -425
rect -1336 -450 -1303 -442
rect -1240 -425 -1207 -417
rect -1240 -442 -1232 -425
rect -1215 -442 -1207 -425
rect -1240 -450 -1207 -442
rect -1144 -424 -1111 -416
rect -1144 -441 -1136 -424
rect -1119 -441 -1111 -424
rect -1144 -449 -1111 -441
rect -1048 -424 -1015 -416
rect -1048 -441 -1040 -424
rect -1023 -441 -1015 -424
rect -1048 -449 -1015 -441
rect -952 -424 -919 -416
rect -952 -441 -944 -424
rect -927 -441 -919 -424
rect -952 -449 -919 -441
rect -856 -424 -823 -416
rect -856 -441 -848 -424
rect -831 -441 -823 -424
rect -856 -449 -823 -441
rect -760 -424 -727 -416
rect -760 -441 -752 -424
rect -735 -441 -727 -424
rect -760 -449 -727 -441
rect -664 -424 -631 -416
rect -664 -441 -656 -424
rect -639 -441 -631 -424
rect -664 -449 -631 -441
rect -568 -424 -535 -416
rect -568 -441 -560 -424
rect -543 -441 -535 -424
rect -568 -449 -535 -441
rect -472 -424 -439 -416
rect -472 -441 -464 -424
rect -447 -441 -439 -424
rect -472 -449 -439 -441
rect -376 -424 -343 -416
rect -376 -441 -368 -424
rect -351 -441 -343 -424
rect -376 -449 -343 -441
rect -280 -424 -247 -416
rect -280 -441 -272 -424
rect -255 -441 -247 -424
rect -280 -449 -247 -441
rect -184 -424 -151 -416
rect -184 -441 -176 -424
rect -159 -441 -151 -424
rect -184 -449 -151 -441
rect -88 -424 -55 -416
rect -88 -441 -80 -424
rect -63 -441 -55 -424
rect -88 -449 -55 -441
rect 7 -424 40 -416
rect 7 -441 15 -424
rect 32 -441 40 -424
rect 7 -449 40 -441
rect 103 -424 136 -416
rect 103 -441 111 -424
rect 128 -441 136 -424
rect 103 -449 136 -441
rect 199 -424 232 -416
rect 199 -441 207 -424
rect 224 -441 232 -424
rect 199 -449 232 -441
rect 295 -424 328 -416
rect 295 -441 303 -424
rect 320 -441 328 -424
rect 295 -449 328 -441
rect 391 -424 424 -416
rect 391 -441 399 -424
rect 416 -441 424 -424
rect 391 -449 424 -441
rect 487 -424 520 -416
rect 487 -441 495 -424
rect 512 -441 520 -424
rect 487 -449 520 -441
rect 583 -424 616 -416
rect 583 -441 591 -424
rect 608 -441 616 -424
rect 583 -449 616 -441
rect 679 -424 712 -416
rect 679 -441 687 -424
rect 704 -441 712 -424
rect 679 -449 712 -441
rect 775 -424 808 -416
rect 775 -441 783 -424
rect 800 -441 808 -424
rect 775 -449 808 -441
rect 871 -424 904 -416
rect 871 -441 879 -424
rect 896 -441 904 -424
rect 871 -449 904 -441
rect 967 -424 1000 -416
rect 967 -441 975 -424
rect 992 -441 1000 -424
rect 967 -449 1000 -441
rect 1063 -424 1096 -416
rect 1063 -441 1071 -424
rect 1088 -441 1096 -424
rect 1063 -449 1096 -441
rect 1159 -424 1192 -416
rect 1159 -441 1167 -424
rect 1184 -441 1192 -424
rect 1159 -449 1192 -441
rect 1255 -424 1288 -416
rect 1255 -441 1263 -424
rect 1280 -441 1288 -424
rect 1255 -449 1288 -441
rect 1351 -424 1384 -416
rect 1351 -441 1359 -424
rect 1376 -441 1384 -424
rect 1351 -449 1384 -441
rect 1447 -424 1480 -416
rect 1447 -441 1455 -424
rect 1472 -441 1480 -424
rect 1447 -449 1480 -441
rect 1543 -424 1576 -416
rect 1543 -441 1551 -424
rect 1568 -441 1576 -424
rect 1543 -449 1576 -441
rect 1639 -424 1672 -416
rect 1639 -441 1647 -424
rect 1664 -441 1672 -424
rect 1639 -449 1672 -441
rect 1735 -424 1768 -416
rect 1735 -441 1743 -424
rect 1760 -441 1768 -424
rect 1735 -449 1768 -441
rect 1831 -424 1864 -416
rect 1831 -441 1839 -424
rect 1856 -441 1864 -424
rect 1831 -449 1864 -441
rect 1927 -424 1960 -416
rect 1927 -441 1935 -424
rect 1952 -441 1960 -424
rect 1927 -449 1960 -441
rect 2023 -424 2056 -416
rect 2023 -441 2031 -424
rect 2048 -441 2056 -424
rect 2023 -449 2056 -441
rect 2119 -424 2152 -416
rect 2119 -441 2127 -424
rect 2144 -441 2152 -424
rect 2119 -449 2152 -441
rect 2215 -424 2248 -416
rect 2215 -441 2223 -424
rect 2240 -441 2248 -424
rect 2215 -449 2248 -441
rect 2311 -424 2344 -416
rect 2311 -441 2319 -424
rect 2336 -441 2344 -424
rect 2311 -449 2344 -441
rect 2407 -424 2440 -416
rect 2407 -441 2415 -424
rect 2432 -441 2440 -424
rect 2407 -449 2440 -441
rect 2503 -424 2536 -416
rect 2503 -441 2511 -424
rect 2528 -441 2536 -424
rect 2503 -449 2536 -441
rect 2599 -424 2632 -416
rect 2599 -441 2607 -424
rect 2624 -441 2632 -424
rect 2599 -449 2632 -441
rect 2695 -424 2728 -416
rect 2695 -441 2703 -424
rect 2720 -441 2728 -424
rect 2695 -449 2728 -441
rect 2791 -424 2824 -416
rect 2791 -441 2799 -424
rect 2816 -441 2824 -424
rect 2791 -449 2824 -441
<< polycont >>
rect -2816 424 -2799 441
rect -2720 424 -2703 441
rect -2624 424 -2607 441
rect -2528 424 -2511 441
rect -2432 424 -2415 441
rect -2336 424 -2319 441
rect -2240 424 -2223 441
rect -2144 424 -2127 441
rect -2048 424 -2031 441
rect -1952 424 -1935 441
rect -1856 424 -1839 441
rect -1760 424 -1743 441
rect -1664 424 -1647 441
rect -1568 424 -1551 441
rect -1472 424 -1455 441
rect -1376 424 -1359 441
rect -1280 424 -1263 441
rect -1184 424 -1167 441
rect -1088 424 -1071 441
rect -992 424 -975 441
rect -896 424 -879 441
rect -800 424 -783 441
rect -704 424 -687 441
rect -608 424 -591 441
rect -512 424 -495 441
rect -416 424 -399 441
rect -320 424 -303 441
rect -224 424 -207 441
rect -128 424 -111 441
rect -32 424 -15 441
rect 63 424 80 441
rect 159 424 176 441
rect 255 424 272 441
rect 351 424 368 441
rect 447 424 464 441
rect 543 424 560 441
rect 639 424 656 441
rect 735 424 752 441
rect 831 424 848 441
rect 927 424 944 441
rect 1023 424 1040 441
rect 1119 424 1136 441
rect 1215 424 1232 441
rect 1311 424 1328 441
rect 1407 424 1424 441
rect 1503 424 1520 441
rect 1599 424 1616 441
rect 1695 424 1712 441
rect 1791 424 1808 441
rect 1887 424 1904 441
rect 1983 424 2000 441
rect 2079 424 2096 441
rect 2175 424 2192 441
rect 2271 424 2288 441
rect 2367 424 2384 441
rect 2463 424 2480 441
rect 2559 424 2576 441
rect 2655 424 2672 441
rect 2751 424 2768 441
rect 2847 424 2864 441
rect -2864 -442 -2847 -425
rect -2768 -442 -2751 -425
rect -2672 -442 -2655 -425
rect -2576 -442 -2559 -425
rect -2480 -442 -2463 -425
rect -2384 -442 -2367 -425
rect -2288 -442 -2271 -425
rect -2192 -442 -2175 -425
rect -2096 -442 -2079 -425
rect -2000 -442 -1983 -425
rect -1904 -442 -1887 -425
rect -1808 -442 -1791 -425
rect -1712 -442 -1695 -425
rect -1616 -442 -1599 -425
rect -1520 -442 -1503 -425
rect -1424 -442 -1407 -425
rect -1328 -442 -1311 -425
rect -1232 -442 -1215 -425
rect -1136 -441 -1119 -424
rect -1040 -441 -1023 -424
rect -944 -441 -927 -424
rect -848 -441 -831 -424
rect -752 -441 -735 -424
rect -656 -441 -639 -424
rect -560 -441 -543 -424
rect -464 -441 -447 -424
rect -368 -441 -351 -424
rect -272 -441 -255 -424
rect -176 -441 -159 -424
rect -80 -441 -63 -424
rect 15 -441 32 -424
rect 111 -441 128 -424
rect 207 -441 224 -424
rect 303 -441 320 -424
rect 399 -441 416 -424
rect 495 -441 512 -424
rect 591 -441 608 -424
rect 687 -441 704 -424
rect 783 -441 800 -424
rect 879 -441 896 -424
rect 975 -441 992 -424
rect 1071 -441 1088 -424
rect 1167 -441 1184 -424
rect 1263 -441 1280 -424
rect 1359 -441 1376 -424
rect 1455 -441 1472 -424
rect 1551 -441 1568 -424
rect 1647 -441 1664 -424
rect 1743 -441 1760 -424
rect 1839 -441 1856 -424
rect 1935 -441 1952 -424
rect 2031 -441 2048 -424
rect 2127 -441 2144 -424
rect 2223 -441 2240 -424
rect 2319 -441 2336 -424
rect 2415 -441 2432 -424
rect 2511 -441 2528 -424
rect 2607 -441 2624 -424
rect 2703 -441 2720 -424
rect 2799 -441 2816 -424
<< locali >>
rect -2945 474 -2897 491
rect 2897 474 2945 491
rect -2945 443 -2928 474
rect 2928 443 2945 474
rect -2824 424 -2816 441
rect -2799 424 -2791 441
rect -2728 424 -2720 441
rect -2703 424 -2695 441
rect -2632 424 -2624 441
rect -2607 424 -2599 441
rect -2536 424 -2528 441
rect -2511 424 -2503 441
rect -2440 424 -2432 441
rect -2415 424 -2407 441
rect -2344 424 -2336 441
rect -2319 424 -2311 441
rect -2248 424 -2240 441
rect -2223 424 -2215 441
rect -2152 424 -2144 441
rect -2127 424 -2119 441
rect -2056 424 -2048 441
rect -2031 424 -2023 441
rect -1960 424 -1952 441
rect -1935 424 -1927 441
rect -1864 424 -1856 441
rect -1839 424 -1831 441
rect -1768 424 -1760 441
rect -1743 424 -1735 441
rect -1672 424 -1664 441
rect -1647 424 -1639 441
rect -1576 424 -1568 441
rect -1551 424 -1543 441
rect -1480 424 -1472 441
rect -1455 424 -1447 441
rect -1384 424 -1376 441
rect -1359 424 -1351 441
rect -1288 424 -1280 441
rect -1263 424 -1255 441
rect -1192 424 -1184 441
rect -1167 424 -1159 441
rect -1096 424 -1088 441
rect -1071 424 -1063 441
rect -1000 424 -992 441
rect -975 424 -967 441
rect -904 424 -896 441
rect -879 424 -871 441
rect -808 424 -800 441
rect -783 424 -775 441
rect -712 424 -704 441
rect -687 424 -679 441
rect -616 424 -608 441
rect -591 424 -583 441
rect -520 424 -512 441
rect -495 424 -487 441
rect -424 424 -416 441
rect -399 424 -391 441
rect -328 424 -320 441
rect -303 424 -295 441
rect -232 424 -224 441
rect -207 424 -199 441
rect -136 424 -128 441
rect -111 424 -103 441
rect -40 424 -32 441
rect -15 424 -7 441
rect 55 424 63 441
rect 80 424 88 441
rect 151 424 159 441
rect 176 424 184 441
rect 247 424 255 441
rect 272 424 280 441
rect 343 424 351 441
rect 368 424 376 441
rect 439 424 447 441
rect 464 424 472 441
rect 535 424 543 441
rect 560 424 568 441
rect 631 424 639 441
rect 656 424 664 441
rect 727 424 735 441
rect 752 424 760 441
rect 823 424 831 441
rect 848 424 856 441
rect 919 424 927 441
rect 944 424 952 441
rect 1015 424 1023 441
rect 1040 424 1048 441
rect 1111 424 1119 441
rect 1136 424 1144 441
rect 1207 424 1215 441
rect 1232 424 1240 441
rect 1303 424 1311 441
rect 1328 424 1336 441
rect 1399 424 1407 441
rect 1424 424 1432 441
rect 1495 424 1503 441
rect 1520 424 1528 441
rect 1591 424 1599 441
rect 1616 424 1624 441
rect 1687 424 1695 441
rect 1712 424 1720 441
rect 1783 424 1791 441
rect 1808 424 1816 441
rect 1879 424 1887 441
rect 1904 424 1912 441
rect 1975 424 1983 441
rect 2000 424 2008 441
rect 2071 424 2079 441
rect 2096 424 2104 441
rect 2167 424 2175 441
rect 2192 424 2200 441
rect 2263 424 2271 441
rect 2288 424 2296 441
rect 2359 424 2367 441
rect 2384 424 2392 441
rect 2455 424 2463 441
rect 2480 424 2488 441
rect 2551 424 2559 441
rect 2576 424 2584 441
rect 2647 424 2655 441
rect 2672 424 2680 441
rect 2743 424 2751 441
rect 2768 424 2776 441
rect 2839 424 2847 441
rect 2864 424 2872 441
rect -2888 394 -2871 402
rect -2888 -402 -2871 -394
rect -2840 394 -2823 402
rect -2840 -402 -2823 -394
rect -2792 394 -2775 402
rect -2792 -402 -2775 -394
rect -2744 394 -2727 402
rect -2744 -402 -2727 -394
rect -2696 394 -2679 402
rect -2696 -402 -2679 -394
rect -2648 394 -2631 402
rect -2648 -402 -2631 -394
rect -2600 394 -2583 402
rect -2600 -402 -2583 -394
rect -2552 394 -2535 402
rect -2552 -402 -2535 -394
rect -2504 394 -2487 402
rect -2504 -402 -2487 -394
rect -2456 394 -2439 402
rect -2456 -402 -2439 -394
rect -2408 394 -2391 402
rect -2408 -402 -2391 -394
rect -2360 394 -2343 402
rect -2360 -402 -2343 -394
rect -2312 394 -2295 402
rect -2312 -402 -2295 -394
rect -2264 394 -2247 402
rect -2264 -402 -2247 -394
rect -2216 394 -2199 402
rect -2216 -402 -2199 -394
rect -2168 394 -2151 402
rect -2168 -402 -2151 -394
rect -2120 394 -2103 402
rect -2120 -402 -2103 -394
rect -2072 394 -2055 402
rect -2072 -402 -2055 -394
rect -2024 394 -2007 402
rect -2024 -402 -2007 -394
rect -1976 394 -1959 402
rect -1976 -402 -1959 -394
rect -1928 394 -1911 402
rect -1928 -402 -1911 -394
rect -1880 394 -1863 402
rect -1880 -402 -1863 -394
rect -1832 394 -1815 402
rect -1832 -402 -1815 -394
rect -1784 394 -1767 402
rect -1784 -402 -1767 -394
rect -1736 394 -1719 402
rect -1736 -402 -1719 -394
rect -1688 394 -1671 402
rect -1688 -402 -1671 -394
rect -1640 394 -1623 402
rect -1640 -402 -1623 -394
rect -1592 394 -1575 402
rect -1592 -402 -1575 -394
rect -1544 394 -1527 402
rect -1544 -402 -1527 -394
rect -1496 394 -1479 402
rect -1496 -402 -1479 -394
rect -1448 394 -1431 402
rect -1448 -402 -1431 -394
rect -1400 394 -1383 402
rect -1400 -402 -1383 -394
rect -1352 394 -1335 402
rect -1352 -402 -1335 -394
rect -1304 394 -1287 402
rect -1304 -402 -1287 -394
rect -1256 394 -1239 402
rect -1256 -402 -1239 -394
rect -1208 394 -1191 402
rect -1208 -402 -1191 -394
rect -1160 394 -1143 402
rect -1160 -402 -1143 -394
rect -1112 394 -1095 402
rect -1112 -402 -1095 -394
rect -1064 394 -1047 402
rect -1064 -402 -1047 -394
rect -1016 394 -999 402
rect -1016 -402 -999 -394
rect -968 394 -951 402
rect -968 -402 -951 -394
rect -920 394 -903 402
rect -920 -402 -903 -394
rect -872 394 -855 402
rect -872 -402 -855 -394
rect -824 394 -807 402
rect -824 -402 -807 -394
rect -776 394 -759 402
rect -776 -402 -759 -394
rect -728 394 -711 402
rect -728 -402 -711 -394
rect -680 394 -663 402
rect -680 -402 -663 -394
rect -632 394 -615 402
rect -632 -402 -615 -394
rect -584 394 -567 402
rect -584 -402 -567 -394
rect -536 394 -519 402
rect -536 -402 -519 -394
rect -488 394 -471 402
rect -488 -402 -471 -394
rect -440 394 -423 402
rect -440 -402 -423 -394
rect -392 394 -375 402
rect -392 -402 -375 -394
rect -344 394 -327 402
rect -344 -402 -327 -394
rect -296 394 -279 402
rect -296 -402 -279 -394
rect -248 394 -231 402
rect -248 -402 -231 -394
rect -200 394 -183 402
rect -200 -402 -183 -394
rect -152 394 -135 402
rect -152 -402 -135 -394
rect -104 394 -87 402
rect -104 -402 -87 -394
rect -56 394 -39 402
rect -56 -402 -39 -394
rect -8 394 9 402
rect -8 -402 9 -394
rect 39 394 56 402
rect 39 -402 56 -394
rect 87 394 104 402
rect 87 -402 104 -394
rect 135 394 152 402
rect 135 -402 152 -394
rect 183 394 200 402
rect 183 -402 200 -394
rect 231 394 248 402
rect 231 -402 248 -394
rect 279 394 296 402
rect 279 -402 296 -394
rect 327 394 344 402
rect 327 -402 344 -394
rect 375 394 392 402
rect 375 -402 392 -394
rect 423 394 440 402
rect 423 -402 440 -394
rect 471 394 488 402
rect 471 -402 488 -394
rect 519 394 536 402
rect 519 -402 536 -394
rect 567 394 584 402
rect 567 -402 584 -394
rect 615 394 632 402
rect 615 -402 632 -394
rect 663 394 680 402
rect 663 -402 680 -394
rect 711 394 728 402
rect 711 -402 728 -394
rect 759 394 776 402
rect 759 -402 776 -394
rect 807 394 824 402
rect 807 -402 824 -394
rect 855 394 872 402
rect 855 -402 872 -394
rect 903 394 920 402
rect 903 -402 920 -394
rect 951 394 968 402
rect 951 -402 968 -394
rect 999 394 1016 402
rect 999 -402 1016 -394
rect 1047 394 1064 402
rect 1047 -402 1064 -394
rect 1095 394 1112 402
rect 1095 -402 1112 -394
rect 1143 394 1160 402
rect 1143 -402 1160 -394
rect 1191 394 1208 402
rect 1191 -402 1208 -394
rect 1239 394 1256 402
rect 1239 -402 1256 -394
rect 1287 394 1304 402
rect 1287 -402 1304 -394
rect 1335 394 1352 402
rect 1335 -402 1352 -394
rect 1383 394 1400 402
rect 1383 -402 1400 -394
rect 1431 394 1448 402
rect 1431 -402 1448 -394
rect 1479 394 1496 402
rect 1479 -402 1496 -394
rect 1527 394 1544 402
rect 1527 -402 1544 -394
rect 1575 394 1592 402
rect 1575 -402 1592 -394
rect 1623 394 1640 402
rect 1623 -402 1640 -394
rect 1671 394 1688 402
rect 1671 -402 1688 -394
rect 1719 394 1736 402
rect 1719 -402 1736 -394
rect 1767 394 1784 402
rect 1767 -402 1784 -394
rect 1815 394 1832 402
rect 1815 -402 1832 -394
rect 1863 394 1880 402
rect 1863 -402 1880 -394
rect 1911 394 1928 402
rect 1911 -402 1928 -394
rect 1959 394 1976 402
rect 1959 -402 1976 -394
rect 2007 394 2024 402
rect 2007 -402 2024 -394
rect 2055 394 2072 402
rect 2055 -402 2072 -394
rect 2103 394 2120 402
rect 2103 -402 2120 -394
rect 2151 394 2168 402
rect 2151 -402 2168 -394
rect 2199 394 2216 402
rect 2199 -402 2216 -394
rect 2247 394 2264 402
rect 2247 -402 2264 -394
rect 2295 394 2312 402
rect 2295 -402 2312 -394
rect 2343 394 2360 402
rect 2343 -402 2360 -394
rect 2391 394 2408 402
rect 2391 -402 2408 -394
rect 2439 394 2456 402
rect 2439 -402 2456 -394
rect 2487 394 2504 402
rect 2487 -402 2504 -394
rect 2535 394 2552 402
rect 2535 -402 2552 -394
rect 2583 394 2600 402
rect 2583 -402 2600 -394
rect 2631 394 2648 402
rect 2631 -402 2648 -394
rect 2679 394 2696 402
rect 2679 -402 2696 -394
rect 2727 394 2744 402
rect 2727 -402 2744 -394
rect 2775 394 2792 402
rect 2775 -402 2792 -394
rect 2823 394 2840 402
rect 2823 -402 2840 -394
rect 2871 394 2888 402
rect 2871 -402 2888 -394
rect -2872 -442 -2864 -425
rect -2847 -442 -2839 -425
rect -2776 -442 -2768 -425
rect -2751 -442 -2743 -425
rect -2680 -442 -2672 -425
rect -2655 -442 -2647 -425
rect -2584 -442 -2576 -425
rect -2559 -442 -2551 -425
rect -2488 -442 -2480 -425
rect -2463 -442 -2455 -425
rect -2392 -442 -2384 -425
rect -2367 -442 -2359 -425
rect -2296 -442 -2288 -425
rect -2271 -442 -2263 -425
rect -2200 -442 -2192 -425
rect -2175 -442 -2167 -425
rect -2104 -442 -2096 -425
rect -2079 -442 -2071 -425
rect -2008 -442 -2000 -425
rect -1983 -442 -1975 -425
rect -1912 -442 -1904 -425
rect -1887 -442 -1879 -425
rect -1816 -442 -1808 -425
rect -1791 -442 -1783 -425
rect -1720 -442 -1712 -425
rect -1695 -442 -1687 -425
rect -1624 -442 -1616 -425
rect -1599 -442 -1591 -425
rect -1528 -442 -1520 -425
rect -1503 -442 -1495 -425
rect -1432 -442 -1424 -425
rect -1407 -442 -1399 -425
rect -1336 -442 -1328 -425
rect -1311 -442 -1303 -425
rect -1240 -442 -1232 -425
rect -1215 -442 -1207 -425
rect -1144 -441 -1136 -424
rect -1119 -441 -1111 -424
rect -1048 -441 -1040 -424
rect -1023 -441 -1015 -424
rect -952 -441 -944 -424
rect -927 -441 -919 -424
rect -856 -441 -848 -424
rect -831 -441 -823 -424
rect -760 -441 -752 -424
rect -735 -441 -727 -424
rect -664 -441 -656 -424
rect -639 -441 -631 -424
rect -568 -441 -560 -424
rect -543 -441 -535 -424
rect -472 -441 -464 -424
rect -447 -441 -439 -424
rect -376 -441 -368 -424
rect -351 -441 -343 -424
rect -280 -441 -272 -424
rect -255 -441 -247 -424
rect -184 -441 -176 -424
rect -159 -441 -151 -424
rect -88 -441 -80 -424
rect -63 -441 -55 -424
rect 7 -441 15 -424
rect 32 -441 40 -424
rect 103 -441 111 -424
rect 128 -441 136 -424
rect 199 -441 207 -424
rect 224 -441 232 -424
rect 295 -441 303 -424
rect 320 -441 328 -424
rect 391 -441 399 -424
rect 416 -441 424 -424
rect 487 -441 495 -424
rect 512 -441 520 -424
rect 583 -441 591 -424
rect 608 -441 616 -424
rect 679 -441 687 -424
rect 704 -441 712 -424
rect 775 -441 783 -424
rect 800 -441 808 -424
rect 871 -441 879 -424
rect 896 -441 904 -424
rect 967 -441 975 -424
rect 992 -441 1000 -424
rect 1063 -441 1071 -424
rect 1088 -441 1096 -424
rect 1159 -441 1167 -424
rect 1184 -441 1192 -424
rect 1255 -441 1263 -424
rect 1280 -441 1288 -424
rect 1351 -441 1359 -424
rect 1376 -441 1384 -424
rect 1447 -441 1455 -424
rect 1472 -441 1480 -424
rect 1543 -441 1551 -424
rect 1568 -441 1576 -424
rect 1639 -441 1647 -424
rect 1664 -441 1672 -424
rect 1735 -441 1743 -424
rect 1760 -441 1768 -424
rect 1831 -441 1839 -424
rect 1856 -441 1864 -424
rect 1927 -441 1935 -424
rect 1952 -441 1960 -424
rect 2023 -441 2031 -424
rect 2048 -441 2056 -424
rect 2119 -441 2127 -424
rect 2144 -441 2152 -424
rect 2215 -441 2223 -424
rect 2240 -441 2248 -424
rect 2311 -441 2319 -424
rect 2336 -441 2344 -424
rect 2407 -441 2415 -424
rect 2432 -441 2440 -424
rect 2503 -441 2511 -424
rect 2528 -441 2536 -424
rect 2599 -441 2607 -424
rect 2624 -441 2632 -424
rect 2695 -441 2703 -424
rect 2720 -441 2728 -424
rect 2791 -441 2799 -424
rect 2816 -441 2824 -424
rect -2945 -474 -2928 -443
rect 2928 -474 2945 -443
rect -2945 -491 -2897 -474
rect 2897 -491 2945 -474
<< viali >>
rect -2816 424 -2799 441
rect -2720 424 -2703 441
rect -2624 424 -2607 441
rect -2528 424 -2511 441
rect -2432 424 -2415 441
rect -2336 424 -2319 441
rect -2240 424 -2223 441
rect -2144 424 -2127 441
rect -2048 424 -2031 441
rect -1952 424 -1935 441
rect -1856 424 -1839 441
rect -1760 424 -1743 441
rect -1664 424 -1647 441
rect -1568 424 -1551 441
rect -1472 424 -1455 441
rect -1376 424 -1359 441
rect -1280 424 -1263 441
rect -1184 424 -1167 441
rect -1088 424 -1071 441
rect -992 424 -975 441
rect -896 424 -879 441
rect -800 424 -783 441
rect -704 424 -687 441
rect -608 424 -591 441
rect -512 424 -495 441
rect -416 424 -399 441
rect -320 424 -303 441
rect -224 424 -207 441
rect -128 424 -111 441
rect -32 424 -15 441
rect 63 424 80 441
rect 159 424 176 441
rect 255 424 272 441
rect 351 424 368 441
rect 447 424 464 441
rect 543 424 560 441
rect 639 424 656 441
rect 735 424 752 441
rect 831 424 848 441
rect 927 424 944 441
rect 1023 424 1040 441
rect 1119 424 1136 441
rect 1215 424 1232 441
rect 1311 424 1328 441
rect 1407 424 1424 441
rect 1503 424 1520 441
rect 1599 424 1616 441
rect 1695 424 1712 441
rect 1791 424 1808 441
rect 1887 424 1904 441
rect 1983 424 2000 441
rect 2079 424 2096 441
rect 2175 424 2192 441
rect 2271 424 2288 441
rect 2367 424 2384 441
rect 2463 424 2480 441
rect 2559 424 2576 441
rect 2655 424 2672 441
rect 2751 424 2768 441
rect 2847 424 2864 441
rect -2888 -394 -2871 394
rect -2840 -394 -2823 394
rect -2792 -394 -2775 394
rect -2744 -394 -2727 394
rect -2696 -394 -2679 394
rect -2648 -394 -2631 394
rect -2600 -394 -2583 394
rect -2552 -394 -2535 394
rect -2504 -394 -2487 394
rect -2456 -394 -2439 394
rect -2408 -394 -2391 394
rect -2360 -394 -2343 394
rect -2312 -394 -2295 394
rect -2264 -394 -2247 394
rect -2216 -394 -2199 394
rect -2168 -394 -2151 394
rect -2120 -394 -2103 394
rect -2072 -394 -2055 394
rect -2024 -394 -2007 394
rect -1976 -394 -1959 394
rect -1928 -394 -1911 394
rect -1880 -394 -1863 394
rect -1832 -394 -1815 394
rect -1784 -394 -1767 394
rect -1736 -394 -1719 394
rect -1688 -394 -1671 394
rect -1640 -394 -1623 394
rect -1592 -394 -1575 394
rect -1544 -394 -1527 394
rect -1496 -394 -1479 394
rect -1448 -394 -1431 394
rect -1400 -394 -1383 394
rect -1352 -394 -1335 394
rect -1304 -394 -1287 394
rect -1256 -394 -1239 394
rect -1208 -394 -1191 394
rect -1160 -394 -1143 394
rect -1112 -394 -1095 394
rect -1064 -394 -1047 394
rect -1016 -394 -999 394
rect -968 -394 -951 394
rect -920 -394 -903 394
rect -872 -394 -855 394
rect -824 -394 -807 394
rect -776 -394 -759 394
rect -728 -394 -711 394
rect -680 -394 -663 394
rect -632 -394 -615 394
rect -584 -394 -567 394
rect -536 -394 -519 394
rect -488 -394 -471 394
rect -440 -394 -423 394
rect -392 -394 -375 394
rect -344 -394 -327 394
rect -296 -394 -279 394
rect -248 -394 -231 394
rect -200 -394 -183 394
rect -152 -394 -135 394
rect -104 -394 -87 394
rect -56 -394 -39 394
rect -8 -394 9 394
rect 39 -394 56 394
rect 87 -394 104 394
rect 135 -394 152 394
rect 183 -394 200 394
rect 231 -394 248 394
rect 279 -394 296 394
rect 327 -394 344 394
rect 375 -394 392 394
rect 423 -394 440 394
rect 471 -394 488 394
rect 519 -394 536 394
rect 567 -394 584 394
rect 615 -394 632 394
rect 663 -394 680 394
rect 711 -394 728 394
rect 759 -394 776 394
rect 807 -394 824 394
rect 855 -394 872 394
rect 903 -394 920 394
rect 951 -394 968 394
rect 999 -394 1016 394
rect 1047 -394 1064 394
rect 1095 -394 1112 394
rect 1143 -394 1160 394
rect 1191 -394 1208 394
rect 1239 -394 1256 394
rect 1287 -394 1304 394
rect 1335 -394 1352 394
rect 1383 -394 1400 394
rect 1431 -394 1448 394
rect 1479 -394 1496 394
rect 1527 -394 1544 394
rect 1575 -394 1592 394
rect 1623 -394 1640 394
rect 1671 -394 1688 394
rect 1719 -394 1736 394
rect 1767 -394 1784 394
rect 1815 -394 1832 394
rect 1863 -394 1880 394
rect 1911 -394 1928 394
rect 1959 -394 1976 394
rect 2007 -394 2024 394
rect 2055 -394 2072 394
rect 2103 -394 2120 394
rect 2151 -394 2168 394
rect 2199 -394 2216 394
rect 2247 -394 2264 394
rect 2295 -394 2312 394
rect 2343 -394 2360 394
rect 2391 -394 2408 394
rect 2439 -394 2456 394
rect 2487 -394 2504 394
rect 2535 -394 2552 394
rect 2583 -394 2600 394
rect 2631 -394 2648 394
rect 2679 -394 2696 394
rect 2727 -394 2744 394
rect 2775 -394 2792 394
rect 2823 -394 2840 394
rect 2871 -394 2888 394
rect -2864 -442 -2847 -425
rect -2768 -442 -2751 -425
rect -2672 -442 -2655 -425
rect -2576 -442 -2559 -425
rect -2480 -442 -2463 -425
rect -2384 -442 -2367 -425
rect -2288 -442 -2271 -425
rect -2192 -442 -2175 -425
rect -2096 -442 -2079 -425
rect -2000 -442 -1983 -425
rect -1904 -442 -1887 -425
rect -1808 -442 -1791 -425
rect -1712 -442 -1695 -425
rect -1616 -442 -1599 -425
rect -1520 -442 -1503 -425
rect -1424 -442 -1407 -425
rect -1328 -442 -1311 -425
rect -1232 -442 -1215 -425
rect -1136 -441 -1119 -424
rect -1040 -441 -1023 -424
rect -944 -441 -927 -424
rect -848 -441 -831 -424
rect -752 -441 -735 -424
rect -656 -441 -639 -424
rect -560 -441 -543 -424
rect -464 -441 -447 -424
rect -368 -441 -351 -424
rect -272 -441 -255 -424
rect -176 -441 -159 -424
rect -80 -441 -63 -424
rect 15 -441 32 -424
rect 111 -441 128 -424
rect 207 -441 224 -424
rect 303 -441 320 -424
rect 399 -441 416 -424
rect 495 -441 512 -424
rect 591 -441 608 -424
rect 687 -441 704 -424
rect 783 -441 800 -424
rect 879 -441 896 -424
rect 975 -441 992 -424
rect 1071 -441 1088 -424
rect 1167 -441 1184 -424
rect 1263 -441 1280 -424
rect 1359 -441 1376 -424
rect 1455 -441 1472 -424
rect 1551 -441 1568 -424
rect 1647 -441 1664 -424
rect 1743 -441 1760 -424
rect 1839 -441 1856 -424
rect 1935 -441 1952 -424
rect 2031 -441 2048 -424
rect 2127 -441 2144 -424
rect 2223 -441 2240 -424
rect 2319 -441 2336 -424
rect 2415 -441 2432 -424
rect 2511 -441 2528 -424
rect 2607 -441 2624 -424
rect 2703 -441 2720 -424
rect 2799 -441 2816 -424
<< metal1 >>
rect -2822 441 -2793 444
rect -2822 424 -2816 441
rect -2799 424 -2793 441
rect -2822 421 -2793 424
rect -2726 441 -2697 444
rect -2726 424 -2720 441
rect -2703 424 -2697 441
rect -2726 421 -2697 424
rect -2630 441 -2601 444
rect -2630 424 -2624 441
rect -2607 424 -2601 441
rect -2630 421 -2601 424
rect -2534 441 -2505 444
rect -2534 424 -2528 441
rect -2511 424 -2505 441
rect -2534 421 -2505 424
rect -2438 441 -2409 444
rect -2438 424 -2432 441
rect -2415 424 -2409 441
rect -2438 421 -2409 424
rect -2342 441 -2313 444
rect -2342 424 -2336 441
rect -2319 424 -2313 441
rect -2342 421 -2313 424
rect -2246 441 -2217 444
rect -2246 424 -2240 441
rect -2223 424 -2217 441
rect -2246 421 -2217 424
rect -2150 441 -2121 444
rect -2150 424 -2144 441
rect -2127 424 -2121 441
rect -2150 421 -2121 424
rect -2054 441 -2025 444
rect -2054 424 -2048 441
rect -2031 424 -2025 441
rect -2054 421 -2025 424
rect -1958 441 -1929 444
rect -1958 424 -1952 441
rect -1935 424 -1929 441
rect -1958 421 -1929 424
rect -1862 441 -1833 444
rect -1862 424 -1856 441
rect -1839 424 -1833 441
rect -1862 421 -1833 424
rect -1766 441 -1737 444
rect -1766 424 -1760 441
rect -1743 424 -1737 441
rect -1766 421 -1737 424
rect -1670 441 -1641 444
rect -1670 424 -1664 441
rect -1647 424 -1641 441
rect -1670 421 -1641 424
rect -1574 441 -1545 444
rect -1574 424 -1568 441
rect -1551 424 -1545 441
rect -1574 421 -1545 424
rect -1478 441 -1449 444
rect -1478 424 -1472 441
rect -1455 424 -1449 441
rect -1478 421 -1449 424
rect -1382 441 -1353 444
rect -1382 424 -1376 441
rect -1359 424 -1353 441
rect -1382 421 -1353 424
rect -1286 441 -1257 444
rect -1286 424 -1280 441
rect -1263 424 -1257 441
rect -1286 421 -1257 424
rect -1190 441 -1161 444
rect -1190 424 -1184 441
rect -1167 424 -1161 441
rect -1190 421 -1161 424
rect -1094 441 -1065 444
rect -1094 424 -1088 441
rect -1071 424 -1065 441
rect -1094 421 -1065 424
rect -998 441 -969 444
rect -998 424 -992 441
rect -975 424 -969 441
rect -998 421 -969 424
rect -902 441 -873 444
rect -902 424 -896 441
rect -879 424 -873 441
rect -902 421 -873 424
rect -806 441 -777 444
rect -806 424 -800 441
rect -783 424 -777 441
rect -806 421 -777 424
rect -710 441 -681 444
rect -710 424 -704 441
rect -687 424 -681 441
rect -710 421 -681 424
rect -614 441 -585 444
rect -614 424 -608 441
rect -591 424 -585 441
rect -614 421 -585 424
rect -518 441 -489 444
rect -518 424 -512 441
rect -495 424 -489 441
rect -518 421 -489 424
rect -422 441 -393 444
rect -422 424 -416 441
rect -399 424 -393 441
rect -422 421 -393 424
rect -326 441 -297 444
rect -326 424 -320 441
rect -303 424 -297 441
rect -326 421 -297 424
rect -230 441 -201 444
rect -230 424 -224 441
rect -207 424 -201 441
rect -230 421 -201 424
rect -134 441 -105 444
rect -134 424 -128 441
rect -111 424 -105 441
rect -134 421 -105 424
rect -38 441 -9 444
rect -38 424 -32 441
rect -15 424 -9 441
rect -38 421 -9 424
rect 57 441 86 444
rect 57 424 63 441
rect 80 424 86 441
rect 57 421 86 424
rect 153 441 182 444
rect 153 424 159 441
rect 176 424 182 441
rect 153 421 182 424
rect 249 441 278 444
rect 249 424 255 441
rect 272 424 278 441
rect 249 421 278 424
rect 345 441 374 444
rect 345 424 351 441
rect 368 424 374 441
rect 345 421 374 424
rect 441 441 470 444
rect 441 424 447 441
rect 464 424 470 441
rect 441 421 470 424
rect 537 441 566 444
rect 537 424 543 441
rect 560 424 566 441
rect 537 421 566 424
rect 633 441 662 444
rect 633 424 639 441
rect 656 424 662 441
rect 633 421 662 424
rect 729 441 758 444
rect 729 424 735 441
rect 752 424 758 441
rect 729 421 758 424
rect 825 441 854 444
rect 825 424 831 441
rect 848 424 854 441
rect 825 421 854 424
rect 921 441 950 444
rect 921 424 927 441
rect 944 424 950 441
rect 921 421 950 424
rect 1017 441 1046 444
rect 1017 424 1023 441
rect 1040 424 1046 441
rect 1017 421 1046 424
rect 1113 441 1142 444
rect 1113 424 1119 441
rect 1136 424 1142 441
rect 1113 421 1142 424
rect 1209 441 1238 444
rect 1209 424 1215 441
rect 1232 424 1238 441
rect 1209 421 1238 424
rect 1305 441 1334 444
rect 1305 424 1311 441
rect 1328 424 1334 441
rect 1305 421 1334 424
rect 1401 441 1430 444
rect 1401 424 1407 441
rect 1424 424 1430 441
rect 1401 421 1430 424
rect 1497 441 1526 444
rect 1497 424 1503 441
rect 1520 424 1526 441
rect 1497 421 1526 424
rect 1593 441 1622 444
rect 1593 424 1599 441
rect 1616 424 1622 441
rect 1593 421 1622 424
rect 1689 441 1718 444
rect 1689 424 1695 441
rect 1712 424 1718 441
rect 1689 421 1718 424
rect 1785 441 1814 444
rect 1785 424 1791 441
rect 1808 424 1814 441
rect 1785 421 1814 424
rect 1881 441 1910 444
rect 1881 424 1887 441
rect 1904 424 1910 441
rect 1881 421 1910 424
rect 1977 441 2006 444
rect 1977 424 1983 441
rect 2000 424 2006 441
rect 1977 421 2006 424
rect 2073 441 2102 444
rect 2073 424 2079 441
rect 2096 424 2102 441
rect 2073 421 2102 424
rect 2169 441 2198 444
rect 2169 424 2175 441
rect 2192 424 2198 441
rect 2169 421 2198 424
rect 2265 441 2294 444
rect 2265 424 2271 441
rect 2288 424 2294 441
rect 2265 421 2294 424
rect 2361 441 2390 444
rect 2361 424 2367 441
rect 2384 424 2390 441
rect 2361 421 2390 424
rect 2457 441 2486 444
rect 2457 424 2463 441
rect 2480 424 2486 441
rect 2457 421 2486 424
rect 2553 441 2582 444
rect 2553 424 2559 441
rect 2576 424 2582 441
rect 2553 421 2582 424
rect 2649 441 2678 444
rect 2649 424 2655 441
rect 2672 424 2678 441
rect 2649 421 2678 424
rect 2745 441 2774 444
rect 2745 424 2751 441
rect 2768 424 2774 441
rect 2745 421 2774 424
rect 2841 441 2870 444
rect 2841 424 2847 441
rect 2864 424 2870 441
rect 2841 421 2870 424
rect -2891 394 -2868 400
rect -2891 -394 -2888 394
rect -2871 -394 -2868 394
rect -2891 -400 -2868 -394
rect -2843 394 -2820 400
rect -2843 -394 -2840 394
rect -2823 -394 -2820 394
rect -2843 -400 -2820 -394
rect -2795 394 -2772 400
rect -2795 -394 -2792 394
rect -2775 -394 -2772 394
rect -2795 -400 -2772 -394
rect -2747 394 -2724 400
rect -2747 -394 -2744 394
rect -2727 -394 -2724 394
rect -2747 -400 -2724 -394
rect -2699 394 -2676 400
rect -2699 -394 -2696 394
rect -2679 -394 -2676 394
rect -2699 -400 -2676 -394
rect -2651 394 -2628 400
rect -2651 -394 -2648 394
rect -2631 -394 -2628 394
rect -2651 -400 -2628 -394
rect -2603 394 -2580 400
rect -2603 -394 -2600 394
rect -2583 -394 -2580 394
rect -2603 -400 -2580 -394
rect -2555 394 -2532 400
rect -2555 -394 -2552 394
rect -2535 -394 -2532 394
rect -2555 -400 -2532 -394
rect -2507 394 -2484 400
rect -2507 -394 -2504 394
rect -2487 -394 -2484 394
rect -2507 -400 -2484 -394
rect -2459 394 -2436 400
rect -2459 -394 -2456 394
rect -2439 -394 -2436 394
rect -2459 -400 -2436 -394
rect -2411 394 -2388 400
rect -2411 -394 -2408 394
rect -2391 -394 -2388 394
rect -2411 -400 -2388 -394
rect -2363 394 -2340 400
rect -2363 -394 -2360 394
rect -2343 -394 -2340 394
rect -2363 -400 -2340 -394
rect -2315 394 -2292 400
rect -2315 -394 -2312 394
rect -2295 -394 -2292 394
rect -2315 -400 -2292 -394
rect -2267 394 -2244 400
rect -2267 -394 -2264 394
rect -2247 -394 -2244 394
rect -2267 -400 -2244 -394
rect -2219 394 -2196 400
rect -2219 -394 -2216 394
rect -2199 -394 -2196 394
rect -2219 -400 -2196 -394
rect -2171 394 -2148 400
rect -2171 -394 -2168 394
rect -2151 -394 -2148 394
rect -2171 -400 -2148 -394
rect -2123 394 -2100 400
rect -2123 -394 -2120 394
rect -2103 -394 -2100 394
rect -2123 -400 -2100 -394
rect -2075 394 -2052 400
rect -2075 -394 -2072 394
rect -2055 -394 -2052 394
rect -2075 -400 -2052 -394
rect -2027 394 -2004 400
rect -2027 -394 -2024 394
rect -2007 -394 -2004 394
rect -2027 -400 -2004 -394
rect -1979 394 -1956 400
rect -1979 -394 -1976 394
rect -1959 -394 -1956 394
rect -1979 -400 -1956 -394
rect -1931 394 -1908 400
rect -1931 -394 -1928 394
rect -1911 -394 -1908 394
rect -1931 -400 -1908 -394
rect -1883 394 -1860 400
rect -1883 -394 -1880 394
rect -1863 -394 -1860 394
rect -1883 -400 -1860 -394
rect -1835 394 -1812 400
rect -1835 -394 -1832 394
rect -1815 -394 -1812 394
rect -1835 -400 -1812 -394
rect -1787 394 -1764 400
rect -1787 -394 -1784 394
rect -1767 -394 -1764 394
rect -1787 -400 -1764 -394
rect -1739 394 -1716 400
rect -1739 -394 -1736 394
rect -1719 -394 -1716 394
rect -1739 -400 -1716 -394
rect -1691 394 -1668 400
rect -1691 -394 -1688 394
rect -1671 -394 -1668 394
rect -1691 -400 -1668 -394
rect -1643 394 -1620 400
rect -1643 -394 -1640 394
rect -1623 -394 -1620 394
rect -1643 -400 -1620 -394
rect -1595 394 -1572 400
rect -1595 -394 -1592 394
rect -1575 -394 -1572 394
rect -1595 -400 -1572 -394
rect -1547 394 -1524 400
rect -1547 -394 -1544 394
rect -1527 -394 -1524 394
rect -1547 -400 -1524 -394
rect -1499 394 -1476 400
rect -1499 -394 -1496 394
rect -1479 -394 -1476 394
rect -1499 -400 -1476 -394
rect -1451 394 -1428 400
rect -1451 -394 -1448 394
rect -1431 -394 -1428 394
rect -1451 -400 -1428 -394
rect -1403 394 -1380 400
rect -1403 -394 -1400 394
rect -1383 -394 -1380 394
rect -1403 -400 -1380 -394
rect -1355 394 -1332 400
rect -1355 -394 -1352 394
rect -1335 -394 -1332 394
rect -1355 -400 -1332 -394
rect -1307 394 -1284 400
rect -1307 -394 -1304 394
rect -1287 -394 -1284 394
rect -1307 -400 -1284 -394
rect -1259 394 -1236 400
rect -1259 -394 -1256 394
rect -1239 -394 -1236 394
rect -1259 -400 -1236 -394
rect -1211 394 -1188 400
rect -1211 -394 -1208 394
rect -1191 -394 -1188 394
rect -1211 -400 -1188 -394
rect -1163 394 -1140 400
rect -1163 -394 -1160 394
rect -1143 -394 -1140 394
rect -1163 -400 -1140 -394
rect -1115 394 -1092 400
rect -1115 -394 -1112 394
rect -1095 -394 -1092 394
rect -1115 -400 -1092 -394
rect -1067 394 -1044 400
rect -1067 -394 -1064 394
rect -1047 -394 -1044 394
rect -1067 -400 -1044 -394
rect -1019 394 -996 400
rect -1019 -394 -1016 394
rect -999 -394 -996 394
rect -1019 -400 -996 -394
rect -971 394 -948 400
rect -971 -394 -968 394
rect -951 -394 -948 394
rect -971 -400 -948 -394
rect -923 394 -900 400
rect -923 -394 -920 394
rect -903 -394 -900 394
rect -923 -400 -900 -394
rect -875 394 -852 400
rect -875 -394 -872 394
rect -855 -394 -852 394
rect -875 -400 -852 -394
rect -827 394 -804 400
rect -827 -394 -824 394
rect -807 -394 -804 394
rect -827 -400 -804 -394
rect -779 394 -756 400
rect -779 -394 -776 394
rect -759 -394 -756 394
rect -779 -400 -756 -394
rect -731 394 -708 400
rect -731 -394 -728 394
rect -711 -394 -708 394
rect -731 -400 -708 -394
rect -683 394 -660 400
rect -683 -394 -680 394
rect -663 -394 -660 394
rect -683 -400 -660 -394
rect -635 394 -612 400
rect -635 -394 -632 394
rect -615 -394 -612 394
rect -635 -400 -612 -394
rect -587 394 -564 400
rect -587 -394 -584 394
rect -567 -394 -564 394
rect -587 -400 -564 -394
rect -539 394 -516 400
rect -539 -394 -536 394
rect -519 -394 -516 394
rect -539 -400 -516 -394
rect -491 394 -468 400
rect -491 -394 -488 394
rect -471 -394 -468 394
rect -491 -400 -468 -394
rect -443 394 -420 400
rect -443 -394 -440 394
rect -423 -394 -420 394
rect -443 -400 -420 -394
rect -395 394 -372 400
rect -395 -394 -392 394
rect -375 -394 -372 394
rect -395 -400 -372 -394
rect -347 394 -324 400
rect -347 -394 -344 394
rect -327 -394 -324 394
rect -347 -400 -324 -394
rect -299 394 -276 400
rect -299 -394 -296 394
rect -279 -394 -276 394
rect -299 -400 -276 -394
rect -251 394 -228 400
rect -251 -394 -248 394
rect -231 -394 -228 394
rect -251 -400 -228 -394
rect -203 394 -180 400
rect -203 -394 -200 394
rect -183 -394 -180 394
rect -203 -400 -180 -394
rect -155 394 -132 400
rect -155 -394 -152 394
rect -135 -394 -132 394
rect -155 -400 -132 -394
rect -107 394 -84 400
rect -107 -394 -104 394
rect -87 -394 -84 394
rect -107 -400 -84 -394
rect -59 394 -36 400
rect -59 -394 -56 394
rect -39 -394 -36 394
rect -59 -400 -36 -394
rect -11 394 12 400
rect -11 -394 -8 394
rect 9 -394 12 394
rect -11 -400 12 -394
rect 36 394 59 400
rect 36 -394 39 394
rect 56 -394 59 394
rect 36 -400 59 -394
rect 84 394 107 400
rect 84 -394 87 394
rect 104 -394 107 394
rect 84 -400 107 -394
rect 132 394 155 400
rect 132 -394 135 394
rect 152 -394 155 394
rect 132 -400 155 -394
rect 180 394 203 400
rect 180 -394 183 394
rect 200 -394 203 394
rect 180 -400 203 -394
rect 228 394 251 400
rect 228 -394 231 394
rect 248 -394 251 394
rect 228 -400 251 -394
rect 276 394 299 400
rect 276 -394 279 394
rect 296 -394 299 394
rect 276 -400 299 -394
rect 324 394 347 400
rect 324 -394 327 394
rect 344 -394 347 394
rect 324 -400 347 -394
rect 372 394 395 400
rect 372 -394 375 394
rect 392 -394 395 394
rect 372 -400 395 -394
rect 420 394 443 400
rect 420 -394 423 394
rect 440 -394 443 394
rect 420 -400 443 -394
rect 468 394 491 400
rect 468 -394 471 394
rect 488 -394 491 394
rect 468 -400 491 -394
rect 516 394 539 400
rect 516 -394 519 394
rect 536 -394 539 394
rect 516 -400 539 -394
rect 564 394 587 400
rect 564 -394 567 394
rect 584 -394 587 394
rect 564 -400 587 -394
rect 612 394 635 400
rect 612 -394 615 394
rect 632 -394 635 394
rect 612 -400 635 -394
rect 660 394 683 400
rect 660 -394 663 394
rect 680 -394 683 394
rect 660 -400 683 -394
rect 708 394 731 400
rect 708 -394 711 394
rect 728 -394 731 394
rect 708 -400 731 -394
rect 756 394 779 400
rect 756 -394 759 394
rect 776 -394 779 394
rect 756 -400 779 -394
rect 804 394 827 400
rect 804 -394 807 394
rect 824 -394 827 394
rect 804 -400 827 -394
rect 852 394 875 400
rect 852 -394 855 394
rect 872 -394 875 394
rect 852 -400 875 -394
rect 900 394 923 400
rect 900 -394 903 394
rect 920 -394 923 394
rect 900 -400 923 -394
rect 948 394 971 400
rect 948 -394 951 394
rect 968 -394 971 394
rect 948 -400 971 -394
rect 996 394 1019 400
rect 996 -394 999 394
rect 1016 -394 1019 394
rect 996 -400 1019 -394
rect 1044 394 1067 400
rect 1044 -394 1047 394
rect 1064 -394 1067 394
rect 1044 -400 1067 -394
rect 1092 394 1115 400
rect 1092 -394 1095 394
rect 1112 -394 1115 394
rect 1092 -400 1115 -394
rect 1140 394 1163 400
rect 1140 -394 1143 394
rect 1160 -394 1163 394
rect 1140 -400 1163 -394
rect 1188 394 1211 400
rect 1188 -394 1191 394
rect 1208 -394 1211 394
rect 1188 -400 1211 -394
rect 1236 394 1259 400
rect 1236 -394 1239 394
rect 1256 -394 1259 394
rect 1236 -400 1259 -394
rect 1284 394 1307 400
rect 1284 -394 1287 394
rect 1304 -394 1307 394
rect 1284 -400 1307 -394
rect 1332 394 1355 400
rect 1332 -394 1335 394
rect 1352 -394 1355 394
rect 1332 -400 1355 -394
rect 1380 394 1403 400
rect 1380 -394 1383 394
rect 1400 -394 1403 394
rect 1380 -400 1403 -394
rect 1428 394 1451 400
rect 1428 -394 1431 394
rect 1448 -394 1451 394
rect 1428 -400 1451 -394
rect 1476 394 1499 400
rect 1476 -394 1479 394
rect 1496 -394 1499 394
rect 1476 -400 1499 -394
rect 1524 394 1547 400
rect 1524 -394 1527 394
rect 1544 -394 1547 394
rect 1524 -400 1547 -394
rect 1572 394 1595 400
rect 1572 -394 1575 394
rect 1592 -394 1595 394
rect 1572 -400 1595 -394
rect 1620 394 1643 400
rect 1620 -394 1623 394
rect 1640 -394 1643 394
rect 1620 -400 1643 -394
rect 1668 394 1691 400
rect 1668 -394 1671 394
rect 1688 -394 1691 394
rect 1668 -400 1691 -394
rect 1716 394 1739 400
rect 1716 -394 1719 394
rect 1736 -394 1739 394
rect 1716 -400 1739 -394
rect 1764 394 1787 400
rect 1764 -394 1767 394
rect 1784 -394 1787 394
rect 1764 -400 1787 -394
rect 1812 394 1835 400
rect 1812 -394 1815 394
rect 1832 -394 1835 394
rect 1812 -400 1835 -394
rect 1860 394 1883 400
rect 1860 -394 1863 394
rect 1880 -394 1883 394
rect 1860 -400 1883 -394
rect 1908 394 1931 400
rect 1908 -394 1911 394
rect 1928 -394 1931 394
rect 1908 -400 1931 -394
rect 1956 394 1979 400
rect 1956 -394 1959 394
rect 1976 -394 1979 394
rect 1956 -400 1979 -394
rect 2004 394 2027 400
rect 2004 -394 2007 394
rect 2024 -394 2027 394
rect 2004 -400 2027 -394
rect 2052 394 2075 400
rect 2052 -394 2055 394
rect 2072 -394 2075 394
rect 2052 -400 2075 -394
rect 2100 394 2123 400
rect 2100 -394 2103 394
rect 2120 -394 2123 394
rect 2100 -400 2123 -394
rect 2148 394 2171 400
rect 2148 -394 2151 394
rect 2168 -394 2171 394
rect 2148 -400 2171 -394
rect 2196 394 2219 400
rect 2196 -394 2199 394
rect 2216 -394 2219 394
rect 2196 -400 2219 -394
rect 2244 394 2267 400
rect 2244 -394 2247 394
rect 2264 -394 2267 394
rect 2244 -400 2267 -394
rect 2292 394 2315 400
rect 2292 -394 2295 394
rect 2312 -394 2315 394
rect 2292 -400 2315 -394
rect 2340 394 2363 400
rect 2340 -394 2343 394
rect 2360 -394 2363 394
rect 2340 -400 2363 -394
rect 2388 394 2411 400
rect 2388 -394 2391 394
rect 2408 -394 2411 394
rect 2388 -400 2411 -394
rect 2436 394 2459 400
rect 2436 -394 2439 394
rect 2456 -394 2459 394
rect 2436 -400 2459 -394
rect 2484 394 2507 400
rect 2484 -394 2487 394
rect 2504 -394 2507 394
rect 2484 -400 2507 -394
rect 2532 394 2555 400
rect 2532 -394 2535 394
rect 2552 -394 2555 394
rect 2532 -400 2555 -394
rect 2580 394 2603 400
rect 2580 -394 2583 394
rect 2600 -394 2603 394
rect 2580 -400 2603 -394
rect 2628 394 2651 400
rect 2628 -394 2631 394
rect 2648 -394 2651 394
rect 2628 -400 2651 -394
rect 2676 394 2699 400
rect 2676 -394 2679 394
rect 2696 -394 2699 394
rect 2676 -400 2699 -394
rect 2724 394 2747 400
rect 2724 -394 2727 394
rect 2744 -394 2747 394
rect 2724 -400 2747 -394
rect 2772 394 2795 400
rect 2772 -394 2775 394
rect 2792 -394 2795 394
rect 2772 -400 2795 -394
rect 2820 394 2843 400
rect 2820 -394 2823 394
rect 2840 -394 2843 394
rect 2820 -400 2843 -394
rect 2868 394 2891 400
rect 2868 -394 2871 394
rect 2888 -394 2891 394
rect 2868 -400 2891 -394
rect -2870 -425 -2841 -422
rect -2870 -442 -2864 -425
rect -2847 -442 -2841 -425
rect -2870 -445 -2841 -442
rect -2774 -425 -2745 -422
rect -2774 -442 -2768 -425
rect -2751 -442 -2745 -425
rect -2774 -445 -2745 -442
rect -2678 -425 -2649 -422
rect -2678 -442 -2672 -425
rect -2655 -442 -2649 -425
rect -2678 -445 -2649 -442
rect -2582 -425 -2553 -422
rect -2582 -442 -2576 -425
rect -2559 -442 -2553 -425
rect -2582 -445 -2553 -442
rect -2486 -425 -2457 -422
rect -2486 -442 -2480 -425
rect -2463 -442 -2457 -425
rect -2486 -445 -2457 -442
rect -2390 -425 -2361 -422
rect -2390 -442 -2384 -425
rect -2367 -442 -2361 -425
rect -2390 -445 -2361 -442
rect -2294 -425 -2265 -422
rect -2294 -442 -2288 -425
rect -2271 -442 -2265 -425
rect -2294 -445 -2265 -442
rect -2198 -425 -2169 -422
rect -2198 -442 -2192 -425
rect -2175 -442 -2169 -425
rect -2198 -445 -2169 -442
rect -2102 -425 -2073 -422
rect -2102 -442 -2096 -425
rect -2079 -442 -2073 -425
rect -2102 -445 -2073 -442
rect -2006 -425 -1977 -422
rect -2006 -442 -2000 -425
rect -1983 -442 -1977 -425
rect -2006 -445 -1977 -442
rect -1910 -425 -1881 -422
rect -1910 -442 -1904 -425
rect -1887 -442 -1881 -425
rect -1910 -445 -1881 -442
rect -1814 -425 -1785 -422
rect -1814 -442 -1808 -425
rect -1791 -442 -1785 -425
rect -1814 -445 -1785 -442
rect -1718 -425 -1689 -422
rect -1718 -442 -1712 -425
rect -1695 -442 -1689 -425
rect -1718 -445 -1689 -442
rect -1622 -425 -1593 -422
rect -1622 -442 -1616 -425
rect -1599 -442 -1593 -425
rect -1622 -445 -1593 -442
rect -1526 -425 -1497 -422
rect -1526 -442 -1520 -425
rect -1503 -442 -1497 -425
rect -1526 -445 -1497 -442
rect -1430 -425 -1401 -422
rect -1430 -442 -1424 -425
rect -1407 -442 -1401 -425
rect -1430 -445 -1401 -442
rect -1334 -425 -1305 -422
rect -1334 -442 -1328 -425
rect -1311 -442 -1305 -425
rect -1334 -445 -1305 -442
rect -1238 -425 -1209 -422
rect -1238 -442 -1232 -425
rect -1215 -442 -1209 -425
rect -1238 -445 -1209 -442
rect -1142 -424 -1113 -421
rect -1142 -441 -1136 -424
rect -1119 -441 -1113 -424
rect -1142 -444 -1113 -441
rect -1046 -424 -1017 -421
rect -1046 -441 -1040 -424
rect -1023 -441 -1017 -424
rect -1046 -444 -1017 -441
rect -950 -424 -921 -421
rect -950 -441 -944 -424
rect -927 -441 -921 -424
rect -950 -444 -921 -441
rect -854 -424 -825 -421
rect -854 -441 -848 -424
rect -831 -441 -825 -424
rect -854 -444 -825 -441
rect -758 -424 -729 -421
rect -758 -441 -752 -424
rect -735 -441 -729 -424
rect -758 -444 -729 -441
rect -662 -424 -633 -421
rect -662 -441 -656 -424
rect -639 -441 -633 -424
rect -662 -444 -633 -441
rect -566 -424 -537 -421
rect -566 -441 -560 -424
rect -543 -441 -537 -424
rect -566 -444 -537 -441
rect -470 -424 -441 -421
rect -470 -441 -464 -424
rect -447 -441 -441 -424
rect -470 -444 -441 -441
rect -374 -424 -345 -421
rect -374 -441 -368 -424
rect -351 -441 -345 -424
rect -374 -444 -345 -441
rect -278 -424 -249 -421
rect -278 -441 -272 -424
rect -255 -441 -249 -424
rect -278 -444 -249 -441
rect -182 -424 -153 -421
rect -182 -441 -176 -424
rect -159 -441 -153 -424
rect -182 -444 -153 -441
rect -86 -424 -57 -421
rect -86 -441 -80 -424
rect -63 -441 -57 -424
rect -86 -444 -57 -441
rect 9 -424 38 -421
rect 9 -441 15 -424
rect 32 -441 38 -424
rect 9 -444 38 -441
rect 105 -424 134 -421
rect 105 -441 111 -424
rect 128 -441 134 -424
rect 105 -444 134 -441
rect 201 -424 230 -421
rect 201 -441 207 -424
rect 224 -441 230 -424
rect 201 -444 230 -441
rect 297 -424 326 -421
rect 297 -441 303 -424
rect 320 -441 326 -424
rect 297 -444 326 -441
rect 393 -424 422 -421
rect 393 -441 399 -424
rect 416 -441 422 -424
rect 393 -444 422 -441
rect 489 -424 518 -421
rect 489 -441 495 -424
rect 512 -441 518 -424
rect 489 -444 518 -441
rect 585 -424 614 -421
rect 585 -441 591 -424
rect 608 -441 614 -424
rect 585 -444 614 -441
rect 681 -424 710 -421
rect 681 -441 687 -424
rect 704 -441 710 -424
rect 681 -444 710 -441
rect 777 -424 806 -421
rect 777 -441 783 -424
rect 800 -441 806 -424
rect 777 -444 806 -441
rect 873 -424 902 -421
rect 873 -441 879 -424
rect 896 -441 902 -424
rect 873 -444 902 -441
rect 969 -424 998 -421
rect 969 -441 975 -424
rect 992 -441 998 -424
rect 969 -444 998 -441
rect 1065 -424 1094 -421
rect 1065 -441 1071 -424
rect 1088 -441 1094 -424
rect 1065 -444 1094 -441
rect 1161 -424 1190 -421
rect 1161 -441 1167 -424
rect 1184 -441 1190 -424
rect 1161 -444 1190 -441
rect 1257 -424 1286 -421
rect 1257 -441 1263 -424
rect 1280 -441 1286 -424
rect 1257 -444 1286 -441
rect 1353 -424 1382 -421
rect 1353 -441 1359 -424
rect 1376 -441 1382 -424
rect 1353 -444 1382 -441
rect 1449 -424 1478 -421
rect 1449 -441 1455 -424
rect 1472 -441 1478 -424
rect 1449 -444 1478 -441
rect 1545 -424 1574 -421
rect 1545 -441 1551 -424
rect 1568 -441 1574 -424
rect 1545 -444 1574 -441
rect 1641 -424 1670 -421
rect 1641 -441 1647 -424
rect 1664 -441 1670 -424
rect 1641 -444 1670 -441
rect 1737 -424 1766 -421
rect 1737 -441 1743 -424
rect 1760 -441 1766 -424
rect 1737 -444 1766 -441
rect 1833 -424 1862 -421
rect 1833 -441 1839 -424
rect 1856 -441 1862 -424
rect 1833 -444 1862 -441
rect 1929 -424 1958 -421
rect 1929 -441 1935 -424
rect 1952 -441 1958 -424
rect 1929 -444 1958 -441
rect 2025 -424 2054 -421
rect 2025 -441 2031 -424
rect 2048 -441 2054 -424
rect 2025 -444 2054 -441
rect 2121 -424 2150 -421
rect 2121 -441 2127 -424
rect 2144 -441 2150 -424
rect 2121 -444 2150 -441
rect 2217 -424 2246 -421
rect 2217 -441 2223 -424
rect 2240 -441 2246 -424
rect 2217 -444 2246 -441
rect 2313 -424 2342 -421
rect 2313 -441 2319 -424
rect 2336 -441 2342 -424
rect 2313 -444 2342 -441
rect 2409 -424 2438 -421
rect 2409 -441 2415 -424
rect 2432 -441 2438 -424
rect 2409 -444 2438 -441
rect 2505 -424 2534 -421
rect 2505 -441 2511 -424
rect 2528 -441 2534 -424
rect 2505 -444 2534 -441
rect 2601 -424 2630 -421
rect 2601 -441 2607 -424
rect 2624 -441 2630 -424
rect 2601 -444 2630 -441
rect 2697 -424 2726 -421
rect 2697 -441 2703 -424
rect 2720 -441 2726 -424
rect 2697 -444 2726 -441
rect 2793 -424 2822 -421
rect 2793 -441 2799 -424
rect 2816 -441 2822 -424
rect 2793 -444 2822 -441
<< properties >>
string FIXED_BBOX -2937 -483 2937 483
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8 l 0.15 m 1 nf 120 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
