magic
tech sky130A
magscale 1 2
timestamp 1697193002
<< error_s >>
rect 132 21802 178 21814
rect 132 21768 138 21802
rect 132 21756 178 21768
rect 1660 21706 1706 21718
rect 1660 21672 1666 21706
rect 1660 21660 1706 21672
rect 132 21610 178 21622
rect 132 21576 138 21610
rect 132 21564 178 21576
rect 1660 21514 1706 21526
rect 1660 21480 1666 21514
rect 1660 21468 1706 21480
rect 132 21418 178 21430
rect 132 21384 138 21418
rect 132 21372 178 21384
rect 1660 21322 1706 21334
rect 1660 21288 1666 21322
rect 1660 21276 1706 21288
rect 132 21226 178 21238
rect 132 21192 138 21226
rect 132 21180 178 21192
rect 1660 21130 1706 21142
rect 1660 21096 1666 21130
rect 1660 21084 1706 21096
rect 132 21034 178 21046
rect 132 21000 138 21034
rect 132 20988 178 21000
rect 1660 20938 1706 20950
rect 1660 20904 1666 20938
rect 1660 20892 1706 20904
rect 132 20842 178 20854
rect 132 20808 138 20842
rect 132 20796 178 20808
rect 1660 20746 1706 20758
rect 1660 20712 1666 20746
rect 1660 20700 1706 20712
rect 132 20650 178 20662
rect 132 20616 138 20650
rect 132 20604 178 20616
rect 1660 20554 1706 20566
rect 1660 20520 1666 20554
rect 1660 20508 1706 20520
rect 132 20458 178 20470
rect 132 20424 138 20458
rect 132 20412 178 20424
rect 1660 20362 1706 20374
rect 1660 20328 1666 20362
rect 1660 20316 1706 20328
rect 132 20266 178 20278
rect 132 20232 138 20266
rect 132 20220 178 20232
rect 1660 20170 1706 20182
rect 1660 20136 1666 20170
rect 1660 20124 1706 20136
rect 132 20074 178 20086
rect 132 20040 138 20074
rect 132 20028 178 20040
rect 1660 19978 1706 19990
rect 1660 19944 1666 19978
rect 1660 19932 1706 19944
rect 132 19882 178 19894
rect 132 19848 138 19882
rect 132 19836 178 19848
rect 1660 19786 1706 19798
rect 1660 19752 1666 19786
rect 1660 19740 1706 19752
rect 132 19690 178 19702
rect 132 19656 138 19690
rect 132 19644 178 19656
rect 1660 19594 1706 19606
rect 1660 19560 1666 19594
rect 1660 19548 1706 19560
rect 132 19498 178 19510
rect 132 19464 138 19498
rect 132 19452 178 19464
rect 1660 19402 1706 19414
rect 1660 19368 1666 19402
rect 1660 19356 1706 19368
rect 132 19306 178 19318
rect 132 19272 138 19306
rect 132 19260 178 19272
rect 1660 19210 1706 19222
rect 1660 19176 1666 19210
rect 1660 19164 1706 19176
rect 132 19114 178 19126
rect 132 19080 138 19114
rect 132 19068 178 19080
rect 1660 19018 1706 19030
rect 1660 18984 1666 19018
rect 1660 18972 1706 18984
rect 132 18922 178 18934
rect 132 18888 138 18922
rect 132 18876 178 18888
rect 1660 18826 1706 18838
rect 1660 18792 1666 18826
rect 1660 18780 1706 18792
rect 132 18730 178 18742
rect 132 18696 138 18730
rect 132 18684 178 18696
rect 1660 18634 1706 18646
rect 1660 18600 1666 18634
rect 1660 18588 1706 18600
rect 132 18538 178 18550
rect 132 18504 138 18538
rect 132 18492 178 18504
rect 1660 18442 1706 18454
rect 1660 18408 1666 18442
rect 1660 18396 1706 18408
rect 132 18346 178 18358
rect 132 18312 138 18346
rect 132 18300 178 18312
rect 1660 18250 1706 18262
rect 1660 18216 1666 18250
rect 1660 18204 1706 18216
rect 132 18154 178 18166
rect 132 18120 138 18154
rect 132 18108 178 18120
rect 1660 18058 1706 18070
rect 1660 18024 1666 18058
rect 1660 18012 1706 18024
rect 132 17962 178 17974
rect 132 17928 138 17962
rect 132 17916 178 17928
rect 1660 17866 1706 17878
rect 1660 17832 1666 17866
rect 1660 17820 1706 17832
rect 132 17770 178 17782
rect 132 17736 138 17770
rect 132 17724 178 17736
rect 1660 17674 1706 17686
rect 1660 17640 1666 17674
rect 1660 17628 1706 17640
rect 132 17578 178 17590
rect 132 17544 138 17578
rect 132 17532 178 17544
rect 1660 17482 1706 17494
rect 1660 17448 1666 17482
rect 1660 17436 1706 17448
rect 132 17386 178 17398
rect 132 17352 138 17386
rect 132 17340 178 17352
rect 1660 17290 1706 17302
rect 1660 17256 1666 17290
rect 1660 17244 1706 17256
rect 132 17194 178 17206
rect 132 17160 138 17194
rect 132 17148 178 17160
rect 1660 17098 1706 17110
rect 1660 17064 1666 17098
rect 1660 17052 1706 17064
rect 132 17002 178 17014
rect 132 16968 138 17002
rect 132 16956 178 16968
rect 1660 16906 1706 16918
rect 1660 16872 1666 16906
rect 1660 16860 1706 16872
rect 132 16810 178 16822
rect 132 16776 138 16810
rect 132 16764 178 16776
rect 1660 16714 1706 16726
rect 1660 16680 1666 16714
rect 1660 16668 1706 16680
rect 132 16618 178 16630
rect 132 16584 138 16618
rect 132 16572 178 16584
rect 1660 16522 1706 16534
rect 1660 16488 1666 16522
rect 1660 16476 1706 16488
rect 132 16426 178 16438
rect 132 16392 138 16426
rect 132 16380 178 16392
rect 1660 16330 1706 16342
rect 1660 16296 1666 16330
rect 1660 16284 1706 16296
rect 132 16234 178 16246
rect 132 16200 138 16234
rect 132 16188 178 16200
rect 1660 16138 1706 16150
rect 1660 16104 1666 16138
rect 1660 16092 1706 16104
rect 132 16042 178 16054
rect 132 16008 138 16042
rect 132 15996 178 16008
rect 1660 15946 1706 15958
rect 1660 15912 1666 15946
rect 1660 15900 1706 15912
rect 132 15850 178 15862
rect 132 15816 138 15850
rect 132 15804 178 15816
rect 1660 15754 1706 15766
rect 1660 15720 1666 15754
rect 1660 15708 1706 15720
rect 132 15658 178 15670
rect 132 15624 138 15658
rect 132 15612 178 15624
rect 1660 15562 1706 15574
rect 1660 15528 1666 15562
rect 1660 15516 1706 15528
rect 132 15466 178 15478
rect 132 15432 138 15466
rect 132 15420 178 15432
rect 1660 15370 1706 15382
rect 1660 15336 1666 15370
rect 1660 15324 1706 15336
rect 132 15274 178 15286
rect 132 15240 138 15274
rect 132 15228 178 15240
rect 1660 15178 1706 15190
rect 1660 15144 1666 15178
rect 1660 15132 1706 15144
rect 132 15082 178 15094
rect 132 15048 138 15082
rect 132 15036 178 15048
rect 1660 14986 1706 14998
rect 1660 14952 1666 14986
rect 1660 14940 1706 14952
rect 132 14890 178 14902
rect 132 14856 138 14890
rect 132 14844 178 14856
rect 1660 14794 1706 14806
rect 1660 14760 1666 14794
rect 1660 14748 1706 14760
rect 132 14698 178 14710
rect 132 14664 138 14698
rect 132 14652 178 14664
rect 1660 14602 1706 14614
rect 1660 14568 1666 14602
rect 1660 14556 1706 14568
rect 132 14506 178 14518
rect 132 14472 138 14506
rect 132 14460 178 14472
rect 1660 14410 1706 14422
rect 1660 14376 1666 14410
rect 1660 14364 1706 14376
rect 132 14314 178 14326
rect 132 14280 138 14314
rect 132 14268 178 14280
rect 1660 14218 1706 14230
rect 1660 14184 1666 14218
rect 1660 14172 1706 14184
rect 132 14122 178 14134
rect 132 14088 138 14122
rect 132 14076 178 14088
rect 1660 14026 1706 14038
rect 1660 13992 1666 14026
rect 1660 13980 1706 13992
rect 132 13930 178 13942
rect 132 13896 138 13930
rect 132 13884 178 13896
rect 1660 13834 1706 13846
rect 1660 13800 1666 13834
rect 1660 13788 1706 13800
rect 132 13738 178 13750
rect 132 13704 138 13738
rect 132 13692 178 13704
rect 1660 13642 1706 13654
rect 1660 13608 1666 13642
rect 1660 13596 1706 13608
rect 132 13546 178 13558
rect 132 13512 138 13546
rect 132 13500 178 13512
rect 1660 13450 1706 13462
rect 1660 13416 1666 13450
rect 1660 13404 1706 13416
rect 132 13354 178 13366
rect 132 13320 138 13354
rect 132 13308 178 13320
rect 1660 13258 1706 13270
rect 1660 13224 1666 13258
rect 1660 13212 1706 13224
rect 132 13162 178 13174
rect 132 13128 138 13162
rect 132 13116 178 13128
rect 1660 13066 1706 13078
rect 1660 13032 1666 13066
rect 1660 13020 1706 13032
rect 132 12970 178 12982
rect 132 12936 138 12970
rect 132 12924 178 12936
rect 1660 12874 1706 12886
rect 1660 12840 1666 12874
rect 1660 12828 1706 12840
rect 132 12778 178 12790
rect 132 12744 138 12778
rect 132 12732 178 12744
rect 1660 12682 1706 12694
rect 1660 12648 1666 12682
rect 1660 12636 1706 12648
rect 132 12586 178 12598
rect 132 12552 138 12586
rect 132 12540 178 12552
rect 1660 12490 1706 12502
rect 1660 12456 1666 12490
rect 1660 12444 1706 12456
rect 132 12394 178 12406
rect 132 12360 138 12394
rect 132 12348 178 12360
rect 1660 12298 1706 12310
rect 1660 12264 1666 12298
rect 1660 12252 1706 12264
rect 132 12202 178 12214
rect 132 12168 138 12202
rect 132 12156 178 12168
rect 1660 12106 1706 12118
rect 1660 12072 1666 12106
rect 1660 12060 1706 12072
rect 132 12010 178 12022
rect 132 11976 138 12010
rect 132 11964 178 11976
rect 1660 11914 1706 11926
rect 1660 11880 1666 11914
rect 1660 11868 1706 11880
rect 132 11818 178 11830
rect 132 11784 138 11818
rect 132 11772 178 11784
rect 1660 11722 1706 11734
rect 1660 11688 1666 11722
rect 1660 11676 1706 11688
rect 132 11626 178 11638
rect 132 11592 138 11626
rect 132 11580 178 11592
rect 1660 11530 1706 11542
rect 1660 11496 1666 11530
rect 1660 11484 1706 11496
rect 132 11434 178 11446
rect 132 11400 138 11434
rect 132 11388 178 11400
rect 1660 11338 1706 11350
rect 1660 11304 1666 11338
rect 1660 11292 1706 11304
rect 132 11242 178 11254
rect 132 11208 138 11242
rect 132 11196 178 11208
rect 1660 11146 1706 11158
rect 1660 11112 1666 11146
rect 1660 11100 1706 11112
rect 132 11050 178 11062
rect 132 11016 138 11050
rect 132 11004 178 11016
rect 1660 10954 1706 10966
rect 1660 10920 1666 10954
rect 1660 10908 1706 10920
rect 132 10858 178 10870
rect 132 10824 138 10858
rect 132 10812 178 10824
rect 1660 10762 1706 10774
rect 1660 10728 1666 10762
rect 1660 10716 1706 10728
rect 132 10666 178 10678
rect 132 10632 138 10666
rect 132 10620 178 10632
rect 1660 10570 1706 10582
rect 1660 10536 1666 10570
rect 1660 10524 1706 10536
rect 132 10474 178 10486
rect 132 10440 138 10474
rect 132 10428 178 10440
rect 1660 10378 1706 10390
rect 1660 10344 1666 10378
rect 1660 10332 1706 10344
rect 132 10282 178 10294
rect 132 10248 138 10282
rect 132 10236 178 10248
rect 1660 10186 1706 10198
rect 1660 10152 1666 10186
rect 1660 10140 1706 10152
rect 132 10090 178 10102
rect 132 10056 138 10090
rect 132 10044 178 10056
rect 1660 9994 1706 10006
rect 1660 9960 1666 9994
rect 1660 9948 1706 9960
rect 132 9898 178 9910
rect 132 9864 138 9898
rect 132 9852 178 9864
rect 1660 9802 1706 9814
rect 1660 9768 1666 9802
rect 1660 9756 1706 9768
rect 132 9706 178 9718
rect 132 9672 138 9706
rect 132 9660 178 9672
rect 1660 9610 1706 9622
rect 1660 9576 1666 9610
rect 1660 9564 1706 9576
rect 132 9514 178 9526
rect 132 9480 138 9514
rect 132 9468 178 9480
rect 1660 9418 1706 9430
rect 1660 9384 1666 9418
rect 1660 9372 1706 9384
rect 132 9322 178 9334
rect 132 9288 138 9322
rect 132 9276 178 9288
rect 1660 9226 1706 9238
rect 1660 9192 1666 9226
rect 1660 9180 1706 9192
rect 132 9130 178 9142
rect 132 9096 138 9130
rect 132 9084 178 9096
rect 1660 9034 1706 9046
rect 1660 9000 1666 9034
rect 1660 8988 1706 9000
rect 132 8938 178 8950
rect 132 8904 138 8938
rect 132 8892 178 8904
rect 1660 8842 1706 8854
rect 1660 8808 1666 8842
rect 1660 8796 1706 8808
rect 132 8746 178 8758
rect 132 8712 138 8746
rect 132 8700 178 8712
rect 1660 8650 1706 8662
rect 1660 8616 1666 8650
rect 1660 8604 1706 8616
rect 132 8554 178 8566
rect 132 8520 138 8554
rect 132 8508 178 8520
rect 1660 8458 1706 8470
rect 1660 8424 1666 8458
rect 1660 8412 1706 8424
rect 132 8362 178 8374
rect 132 8328 138 8362
rect 132 8316 178 8328
rect 1660 8266 1706 8278
rect 1660 8232 1666 8266
rect 1660 8220 1706 8232
rect 132 8170 178 8182
rect 132 8136 138 8170
rect 132 8124 178 8136
rect 1660 8074 1706 8086
rect 1660 8040 1666 8074
rect 1660 8028 1706 8040
rect 132 7978 178 7990
rect 132 7944 138 7978
rect 132 7932 178 7944
rect 1660 7882 1706 7894
rect 1660 7848 1666 7882
rect 1660 7836 1706 7848
rect 132 7786 178 7798
rect 132 7752 138 7786
rect 132 7740 178 7752
rect 1660 7690 1706 7702
rect 1660 7656 1666 7690
rect 1660 7644 1706 7656
rect 132 7594 178 7606
rect 132 7560 138 7594
rect 132 7548 178 7560
rect 1660 7498 1706 7510
rect 1660 7464 1666 7498
rect 1660 7452 1706 7464
rect 132 7402 178 7414
rect 132 7368 138 7402
rect 132 7356 178 7368
rect 1660 7306 1706 7318
rect 1660 7272 1666 7306
rect 1660 7260 1706 7272
rect 132 7210 178 7222
rect 132 7176 138 7210
rect 132 7164 178 7176
rect 1660 7114 1706 7126
rect 1660 7080 1666 7114
rect 1660 7068 1706 7080
rect 132 7018 178 7030
rect 132 6984 138 7018
rect 132 6972 178 6984
rect 1660 6922 1706 6934
rect 1660 6888 1666 6922
rect 1660 6876 1706 6888
rect 132 6826 178 6838
rect 132 6792 138 6826
rect 132 6780 178 6792
rect 1660 6730 1706 6742
rect 1660 6696 1666 6730
rect 1660 6684 1706 6696
rect 132 6634 178 6646
rect 132 6600 138 6634
rect 132 6588 178 6600
rect 1660 6538 1706 6550
rect 1660 6504 1666 6538
rect 1660 6492 1706 6504
rect 132 6442 178 6454
rect 132 6408 138 6442
rect 132 6396 178 6408
rect 1660 6346 1706 6358
rect 1660 6312 1666 6346
rect 1660 6300 1706 6312
rect 132 6250 178 6262
rect 132 6216 138 6250
rect 132 6204 178 6216
rect 1660 6154 1706 6166
rect 1660 6120 1666 6154
rect 1660 6108 1706 6120
rect 132 6058 178 6070
rect 132 6024 138 6058
rect 132 6012 178 6024
rect 1660 5962 1706 5974
rect 1660 5928 1666 5962
rect 1660 5916 1706 5928
rect 132 5866 178 5878
rect 132 5832 138 5866
rect 132 5820 178 5832
rect 1660 5770 1706 5782
rect 1660 5736 1666 5770
rect 1660 5724 1706 5736
rect 132 5674 178 5686
rect 132 5640 138 5674
rect 132 5628 178 5640
rect 1660 5578 1706 5590
rect 1660 5544 1666 5578
rect 1660 5532 1706 5544
rect 132 5482 178 5494
rect 132 5448 138 5482
rect 132 5436 178 5448
rect 1660 5386 1706 5398
rect 1660 5352 1666 5386
rect 1660 5340 1706 5352
rect 132 5290 178 5302
rect 132 5256 138 5290
rect 132 5244 178 5256
rect 1660 5194 1706 5206
rect 1660 5160 1666 5194
rect 1660 5148 1706 5160
rect 132 5098 178 5110
rect 132 5064 138 5098
rect 132 5052 178 5064
rect 1660 5002 1706 5014
rect 1660 4968 1666 5002
rect 1660 4956 1706 4968
rect 132 4906 178 4918
rect 132 4872 138 4906
rect 132 4860 178 4872
rect 1660 4810 1706 4822
rect 1660 4776 1666 4810
rect 1660 4764 1706 4776
rect 132 4714 178 4726
rect 132 4680 138 4714
rect 132 4668 178 4680
rect 1660 4618 1706 4630
rect 1660 4584 1666 4618
rect 1660 4572 1706 4584
rect 132 4522 178 4534
rect 132 4488 138 4522
rect 132 4476 178 4488
rect 1660 4426 1706 4438
rect 1660 4392 1666 4426
rect 1660 4380 1706 4392
rect 132 4330 178 4342
rect 132 4296 138 4330
rect 132 4284 178 4296
rect 1660 4234 1706 4246
rect 1660 4200 1666 4234
rect 1660 4188 1706 4200
rect 132 4138 178 4150
rect 132 4104 138 4138
rect 132 4092 178 4104
rect 1660 4042 1706 4054
rect 1660 4008 1666 4042
rect 1660 3996 1706 4008
rect 132 3946 178 3958
rect 132 3912 138 3946
rect 132 3900 178 3912
rect 1660 3850 1706 3862
rect 1660 3816 1666 3850
rect 1660 3804 1706 3816
rect 132 3754 178 3766
rect 132 3720 138 3754
rect 132 3708 178 3720
rect 1660 3658 1706 3670
rect 1660 3624 1666 3658
rect 1660 3612 1706 3624
rect 132 3562 178 3574
rect 132 3528 138 3562
rect 132 3516 178 3528
rect 1660 3466 1706 3478
rect 1660 3432 1666 3466
rect 1660 3420 1706 3432
rect 132 3370 178 3382
rect 132 3336 138 3370
rect 132 3324 178 3336
rect 1660 3274 1706 3286
rect 1660 3240 1666 3274
rect 1660 3228 1706 3240
rect 132 3178 178 3190
rect 132 3144 138 3178
rect 132 3132 178 3144
rect 1660 3082 1706 3094
rect 1660 3048 1666 3082
rect 1660 3036 1706 3048
rect 132 2986 178 2998
rect 132 2952 138 2986
rect 132 2940 178 2952
rect 1660 2890 1706 2902
rect 1660 2856 1666 2890
rect 1660 2844 1706 2856
rect 132 2794 178 2806
rect 132 2760 138 2794
rect 132 2748 178 2760
rect 1660 2698 1706 2710
rect 1660 2664 1666 2698
rect 1660 2652 1706 2664
rect 132 2602 178 2614
rect 132 2568 138 2602
rect 132 2556 178 2568
rect 1660 2506 1706 2518
rect 1660 2472 1666 2506
rect 1660 2460 1706 2472
rect 132 2410 178 2422
rect 132 2376 138 2410
rect 132 2364 178 2376
rect 1660 2314 1706 2326
rect 1660 2280 1666 2314
rect 1660 2268 1706 2280
rect 132 2218 178 2230
rect 132 2184 138 2218
rect 132 2172 178 2184
rect 1660 2122 1706 2134
rect 1660 2088 1666 2122
rect 1660 2076 1706 2088
rect 132 2026 178 2038
rect 132 1992 138 2026
rect 132 1980 178 1992
rect 1660 1930 1706 1942
rect 1660 1896 1666 1930
rect 1660 1884 1706 1896
rect 132 1834 178 1846
rect 132 1800 138 1834
rect 132 1788 178 1800
rect 1660 1738 1706 1750
rect 1660 1704 1666 1738
rect 1660 1692 1706 1704
rect 132 1642 178 1654
rect 132 1608 138 1642
rect 132 1596 178 1608
rect 1660 1546 1706 1558
rect 1660 1512 1666 1546
rect 1660 1500 1706 1512
rect 132 1450 178 1462
rect 132 1416 138 1450
rect 132 1404 178 1416
rect 1660 1354 1706 1366
rect 1660 1320 1666 1354
rect 1660 1308 1706 1320
rect 132 1258 178 1270
rect 132 1224 138 1258
rect 132 1212 178 1224
rect 1660 1162 1706 1174
rect 1660 1128 1666 1162
rect 1660 1116 1706 1128
rect 132 1066 178 1078
rect 132 1032 138 1066
rect 132 1020 178 1032
rect 1660 970 1706 982
rect 1660 936 1666 970
rect 1660 924 1706 936
rect 132 874 178 886
rect 132 840 138 874
rect 132 828 178 840
rect 1660 778 1706 790
rect 1660 744 1666 778
rect 1660 732 1706 744
<< metal4 >>
rect 0 22204 1840 22304
rect 0 0 240 22000
rect 340 0 870 22000
rect 970 0 1500 22000
rect 1600 0 1840 22000
use sky130_fd_pr__pfet_01v8_6QHARF  sky130_fd_pr__pfet_01v8_6QHARF_0
timestamp 1697193002
transform 0 1 919 -1 0 11273
box -10727 -919 10727 919
<< labels >>
rlabel metal4 0 0 240 22000 1 VGND
port 1 n ground input
rlabel metal4 1600 0 1840 22000 1 VGND
port 1 n ground input
rlabel metal4 340 0 870 22000 1 VPWR
port 2 n power input
rlabel metal4 970 0 1500 22000 1 GPWR
port 3 n power output
rlabel metal4 0 22204 1840 22304 1 ctrl
port 4 n signal input
<< end >>
